module top ( 
    A0 , A1 , A2 , A3 , A4 , A5 , A6 , A7 , A8 ,
    A9 , A10 , A11 , A12 , A13 , A14 , A15 , A16 ,
    A17 , A18 , A19 , A20 , A21 , A22 , A23 , A24 ,
    A25 , A26 , A27 , A28 , A29 , A30 , A31 , A32 ,
    A33 , A34 , A35 , A36 , A37 , A38 , A39 , A40 ,
    A41 , A42 , A43 , A44 , A45 , A46 , A47 , A48 ,
    A49 , A50 , A51 , A52 , A53 , A54 , A55 , A56 ,
    A57 , A58 , A59 , A60 , A61 , A62 , A63 , A64 ,
    A65 , A66 , A67 , A68 , A69 , A70 , A71 , A72 ,
    A73 , A74 , A75 , A76 , A77 , A78 , A79 , A80 ,
    A81 , A82 , A83 , A84 , A85 , A86 , A87 , A88 ,
    A89 , A90 , A91 , A92 , A93 , A94 , A95 , A96 ,
    A97 , A98 , A99 , A100 , A101 , A102 , A103 ,
    A104 , A105 , A106 , A107 , A108 , A109 , A110 ,
    A111 , A112 , A113 , A114 , A115 , A116 , A117 ,
    A118 , A119 , A120 , A121 , A122 , A123 , A124 ,
    A125 , A126 , A127 , A128 , A129 , A130 , A131 ,
    A132 , A133 , A134 , A135 , A136 , A137 , A138 ,
    A139 , A140 , A141 , A142 , A143 , A144 , A145 ,
    A146 , A147 , A148 , A149 , A150 , A151 , A152 ,
    A153 , A154 , A155 , A156 , A157 , A158 , A159 ,
    A160 , A161 , A162 , A163 , A164 , A165 , A166 ,
    A167 , A168 , A169 , A170 , A171 , A172 , A173 ,
    A174 , A175 , A176 , A177 , A178 , A179 , A180 ,
    A181 , A182 , A183 , A184 , A185 , A186 , A187 ,
    A188 , A189 , A190 , A191 , A192 , A193 , A194 ,
    A195 , A196 , A197 , A198 , A199 , A200 , A201 ,
    A202 , A203 , A204 , A205 , A206 , A207 , A208 ,
    A209 , A210 , A211 , A212 , A213 , A214 , A215 ,
    A216 , A217 , A218 , A219 , A220 , A221 , A222 ,
    A223 , A224 , A225 , A226 , A227 , A228 , A229 ,
    A230 , A231 , A232 , A233 , A234 , A235 , A236 ,
    A237 , A238 , A239 , A240 , A241 , A242 , A243 ,
    A244 , A245 , A246 , A247 , A248 , A249 , A250 ,
    A251 , A252 , A253 , A254 , A255 , A256 , A257 ,
    A258 , A259 , A260 , A261 , A262 , A263 , A264 ,
    A265 , A266 , A267 , A268 , A269 , A270 , A271 ,
    A272 , A273 , A274 , A275 , A276 , A277 , A278 ,
    A279 , A280 , A281 , A282 , A283 , A284 , A285 ,
    A286 , A287 , A288 , A289 , A290 , A291 , A292 ,
    A293 , A294 , A295 , A296 , A297 , A298 , A299 ,
    A300 , A301 , A302 , A303 , A304 , A305 , A306 ,
    A307 , A308 , A309 , A310 , A311 , A312 , A313 ,
    A314 , A315 , A316 , A317 , A318 , A319 , A320 ,
    A321 , A322 , A323 , A324 , A325 , A326 , A327 ,
    A328 , A329 , A330 , A331 , A332 , A333 , A334 ,
    A335 , A336 , A337 , A338 , A339 , A340 , A341 ,
    A342 , A343 , A344 , A345 , A346 , A347 , A348 ,
    A349 , A350 , A351 , A352 , A353 , A354 , A355 ,
    A356 , A357 , A358 , A359 , A360 , A361 , A362 ,
    A363 , A364 , A365 , A366 , A367 , A368 , A369 ,
    A370 , A371 , A372 , A373 , A374 , A375 , A376 ,
    A377 , A378 , A379 , A380 , A381 , A382 , A383 ,
    A384 , A385 , A386 , A387 , A388 , A389 , A390 ,
    A391 , A392 , A393 , A394 , A395 , A396 , A397 ,
    A398 , A399 , A400 , A401 , A402 , A403 , A404 ,
    A405 , A406 , A407 , A408 , A409 , A410 , A411 ,
    A412 , A413 , A414 , A415 , A416 , A417 , A418 ,
    A419 , A420 , A421 , A422 , A423 , A424 , A425 ,
    A426 , A427 , A428 , A429 , A430 , A431 , A432 ,
    A433 , A434 , A435 , A436 , A437 , A438 , A439 ,
    A440 , A441 , A442 , A443 , A444 , A445 , A446 ,
    A447 , A448 , A449 , A450 , A451 , A452 , A453 ,
    A454 , A455 , A456 , A457 , A458 , A459 , A460 ,
    A461 , A462 , A463 , A464 , A465 , A466 , A467 ,
    A468 , A469 , A470 , A471 , A472 , A473 , A474 ,
    A475 , A476 , A477 , A478 , A479 , A480 , A481 ,
    A482 , A483 , A484 , A485 , A486 , A487 , A488 ,
    A489 , A490 , A491 , A492 , A493 , A494 , A495 ,
    A496 , A497 , A498 , A499 , A500 , A501 , A502 ,
    A503 , A504 , A505 , A506 , A507 , A508 , A509 ,
    A510 , A511 , A512 , A513 , A514 , A515 , A516 ,
    A517 , A518 , A519 , A520 , A521 , A522 , A523 ,
    A524 , A525 , A526 , A527 , A528 , A529 , A530 ,
    A531 , A532 , A533 , A534 , A535 , A536 , A537 ,
    A538 , A539 , A540 , A541 , A542 , A543 , A544 ,
    A545 , A546 , A547 , A548 , A549 , A550 , A551 ,
    A552 , A553 , A554 , A555 , A556 , A557 , A558 ,
    A559 , A560 , A561 , A562 , A563 , A564 , A565 ,
    A566 , A567 , A568 , A569 , A570 , A571 , A572 ,
    A573 , A574 , A575 , A576 , A577 , A578 , A579 ,
    A580 , A581 , A582 , A583 , A584 , A585 , A586 ,
    A587 , A588 , A589 , A590 , A591 , A592 , A593 ,
    A594 , A595 , A596 , A597 , A598 , A599 , A600 ,
    A601 , A602 , A603 , A604 , A605 , A606 , A607 ,
    A608 , A609 , A610 , A611 , A612 , A613 , A614 ,
    A615 , A616 , A617 , A618 , A619 , A620 , A621 ,
    A622 , A623 , A624 , A625 , A626 , A627 , A628 ,
    A629 , A630 , A631 , A632 , A633 , A634 , A635 ,
    A636 , A637 , A638 , A639 , A640 , A641 , A642 ,
    A643 , A644 , A645 , A646 , A647 , A648 , A649 ,
    A650 , A651 , A652 , A653 , A654 , A655 , A656 ,
    A657 , A658 , A659 , A660 , A661 , A662 , A663 ,
    A664 , A665 , A666 , A667 , A668 , A669 , A670 ,
    A671 , A672 , A673 , A674 , A675 , A676 , A677 ,
    A678 , A679 , A680 , A681 , A682 , A683 , A684 ,
    A685 , A686 , A687 , A688 , A689 , A690 , A691 ,
    A692 , A693 , A694 , A695 , A696 , A697 , A698 ,
    A699 , A700 , A701 , A702 , A703 , A704 , A705 ,
    A706 , A707 , A708 , A709 , A710 , A711 , A712 ,
    A713 , A714 , A715 , A716 , A717 , A718 , A719 ,
    A720 , A721 , A722 , A723 , A724 , A725 , A726 ,
    A727 , A728 , A729 , A730 , A731 , A732 , A733 ,
    A734 , A735 , A736 , A737 , A738 , A739 , A740 ,
    A741 , A742 , A743 , A744 , A745 , A746 , A747 ,
    A748 , A749 , A750 , A751 , A752 , A753 , A754 ,
    A755 , A756 , A757 , A758 , A759 , A760 , A761 ,
    A762 , A763 , A764 , A765 , A766 , A767 , A768 ,
    A769 , A770 , A771 , A772 , A773 , A774 , A775 ,
    A776 , A777 , A778 , A779 , A780 , A781 , A782 ,
    A783 , A784 , A785 , A786 , A787 , A788 , A789 ,
    A790 , A791 , A792 , A793 , A794 , A795 , A796 ,
    A797 , A798 , A799 , A800 , A801 , A802 , A803 ,
    A804 , A805 , A806 , A807 , A808 , A809 , A810 ,
    A811 , A812 , A813 , A814 , A815 , A816 , A817 ,
    A818 , A819 , A820 , A821 , A822 , A823 , A824 ,
    A825 , A826 , A827 , A828 , A829 , A830 , A831 ,
    A832 , A833 , A834 , A835 , A836 , A837 , A838 ,
    A839 , A840 , A841 , A842 , A843 , A844 , A845 ,
    A846 , A847 , A848 , A849 , A850 , A851 , A852 ,
    A853 , A854 , A855 , A856 , A857 , A858 , A859 ,
    A860 , A861 , A862 , A863 , A864 , A865 , A866 ,
    A867 , A868 , A869 , A870 , A871 , A872 , A873 ,
    A874 , A875 , A876 , A877 , A878 , A879 , A880 ,
    A881 , A882 , A883 , A884 , A885 , A886 , A887 ,
    A888 , A889 , A890 , A891 , A892 , A893 , A894 ,
    A895 , A896 , A897 , A898 , A899 , A900 , A901 ,
    A902 , A903 , A904 , A905 , A906 , A907 , A908 ,
    A909 , A910 , A911 , A912 , A913 , A914 , A915 ,
    A916 , A917 , A918 , A919 , A920 , A921 , A922 ,
    A923 , A924 , A925 , A926 , A927 , A928 , A929 ,
    A930 , A931 , A932 , A933 , A934 , A935 , A936 ,
    A937 , A938 , A939 , A940 , A941 , A942 , A943 ,
    A944 , A945 , A946 , A947 , A948 , A949 , A950 ,
    A951 , A952 , A953 , A954 , A955 , A956 , A957 ,
    A958 , A959 , A960 , A961 , A962 , A963 , A964 ,
    A965 , A966 , A967 , A968 , A969 , A970 , A971 ,
    A972 , A973 , A974 , A975 , A976 , A977 , A978 ,
    A979 , A980 , A981 , A982 , A983 , A984 , A985 ,
    A986 , A987 , A988 , A989 , A990 , A991 , A992 ,
    A993 , A994 , A995 , A996 , A997 , A998 , A999 ,
    A1000 ,
    maj  );
  input  A0 , A1 , A2 , A3 , A4 , A5 , A6 , A7 ,
    A8 , A9 , A10 , A11 , A12 , A13 , A14 , A15 ,
    A16 , A17 , A18 , A19 , A20 , A21 , A22 , A23 ,
    A24 , A25 , A26 , A27 , A28 , A29 , A30 , A31 ,
    A32 , A33 , A34 , A35 , A36 , A37 , A38 , A39 ,
    A40 , A41 , A42 , A43 , A44 , A45 , A46 , A47 ,
    A48 , A49 , A50 , A51 , A52 , A53 , A54 , A55 ,
    A56 , A57 , A58 , A59 , A60 , A61 , A62 , A63 ,
    A64 , A65 , A66 , A67 , A68 , A69 , A70 , A71 ,
    A72 , A73 , A74 , A75 , A76 , A77 , A78 , A79 ,
    A80 , A81 , A82 , A83 , A84 , A85 , A86 , A87 ,
    A88 , A89 , A90 , A91 , A92 , A93 , A94 , A95 ,
    A96 , A97 , A98 , A99 , A100 , A101 , A102 ,
    A103 , A104 , A105 , A106 , A107 , A108 , A109 ,
    A110 , A111 , A112 , A113 , A114 , A115 , A116 ,
    A117 , A118 , A119 , A120 , A121 , A122 , A123 ,
    A124 , A125 , A126 , A127 , A128 , A129 , A130 ,
    A131 , A132 , A133 , A134 , A135 , A136 , A137 ,
    A138 , A139 , A140 , A141 , A142 , A143 , A144 ,
    A145 , A146 , A147 , A148 , A149 , A150 , A151 ,
    A152 , A153 , A154 , A155 , A156 , A157 , A158 ,
    A159 , A160 , A161 , A162 , A163 , A164 , A165 ,
    A166 , A167 , A168 , A169 , A170 , A171 , A172 ,
    A173 , A174 , A175 , A176 , A177 , A178 , A179 ,
    A180 , A181 , A182 , A183 , A184 , A185 , A186 ,
    A187 , A188 , A189 , A190 , A191 , A192 , A193 ,
    A194 , A195 , A196 , A197 , A198 , A199 , A200 ,
    A201 , A202 , A203 , A204 , A205 , A206 , A207 ,
    A208 , A209 , A210 , A211 , A212 , A213 , A214 ,
    A215 , A216 , A217 , A218 , A219 , A220 , A221 ,
    A222 , A223 , A224 , A225 , A226 , A227 , A228 ,
    A229 , A230 , A231 , A232 , A233 , A234 , A235 ,
    A236 , A237 , A238 , A239 , A240 , A241 , A242 ,
    A243 , A244 , A245 , A246 , A247 , A248 , A249 ,
    A250 , A251 , A252 , A253 , A254 , A255 , A256 ,
    A257 , A258 , A259 , A260 , A261 , A262 , A263 ,
    A264 , A265 , A266 , A267 , A268 , A269 , A270 ,
    A271 , A272 , A273 , A274 , A275 , A276 , A277 ,
    A278 , A279 , A280 , A281 , A282 , A283 , A284 ,
    A285 , A286 , A287 , A288 , A289 , A290 , A291 ,
    A292 , A293 , A294 , A295 , A296 , A297 , A298 ,
    A299 , A300 , A301 , A302 , A303 , A304 , A305 ,
    A306 , A307 , A308 , A309 , A310 , A311 , A312 ,
    A313 , A314 , A315 , A316 , A317 , A318 , A319 ,
    A320 , A321 , A322 , A323 , A324 , A325 , A326 ,
    A327 , A328 , A329 , A330 , A331 , A332 , A333 ,
    A334 , A335 , A336 , A337 , A338 , A339 , A340 ,
    A341 , A342 , A343 , A344 , A345 , A346 , A347 ,
    A348 , A349 , A350 , A351 , A352 , A353 , A354 ,
    A355 , A356 , A357 , A358 , A359 , A360 , A361 ,
    A362 , A363 , A364 , A365 , A366 , A367 , A368 ,
    A369 , A370 , A371 , A372 , A373 , A374 , A375 ,
    A376 , A377 , A378 , A379 , A380 , A381 , A382 ,
    A383 , A384 , A385 , A386 , A387 , A388 , A389 ,
    A390 , A391 , A392 , A393 , A394 , A395 , A396 ,
    A397 , A398 , A399 , A400 , A401 , A402 , A403 ,
    A404 , A405 , A406 , A407 , A408 , A409 , A410 ,
    A411 , A412 , A413 , A414 , A415 , A416 , A417 ,
    A418 , A419 , A420 , A421 , A422 , A423 , A424 ,
    A425 , A426 , A427 , A428 , A429 , A430 , A431 ,
    A432 , A433 , A434 , A435 , A436 , A437 , A438 ,
    A439 , A440 , A441 , A442 , A443 , A444 , A445 ,
    A446 , A447 , A448 , A449 , A450 , A451 , A452 ,
    A453 , A454 , A455 , A456 , A457 , A458 , A459 ,
    A460 , A461 , A462 , A463 , A464 , A465 , A466 ,
    A467 , A468 , A469 , A470 , A471 , A472 , A473 ,
    A474 , A475 , A476 , A477 , A478 , A479 , A480 ,
    A481 , A482 , A483 , A484 , A485 , A486 , A487 ,
    A488 , A489 , A490 , A491 , A492 , A493 , A494 ,
    A495 , A496 , A497 , A498 , A499 , A500 , A501 ,
    A502 , A503 , A504 , A505 , A506 , A507 , A508 ,
    A509 , A510 , A511 , A512 , A513 , A514 , A515 ,
    A516 , A517 , A518 , A519 , A520 , A521 , A522 ,
    A523 , A524 , A525 , A526 , A527 , A528 , A529 ,
    A530 , A531 , A532 , A533 , A534 , A535 , A536 ,
    A537 , A538 , A539 , A540 , A541 , A542 , A543 ,
    A544 , A545 , A546 , A547 , A548 , A549 , A550 ,
    A551 , A552 , A553 , A554 , A555 , A556 , A557 ,
    A558 , A559 , A560 , A561 , A562 , A563 , A564 ,
    A565 , A566 , A567 , A568 , A569 , A570 , A571 ,
    A572 , A573 , A574 , A575 , A576 , A577 , A578 ,
    A579 , A580 , A581 , A582 , A583 , A584 , A585 ,
    A586 , A587 , A588 , A589 , A590 , A591 , A592 ,
    A593 , A594 , A595 , A596 , A597 , A598 , A599 ,
    A600 , A601 , A602 , A603 , A604 , A605 , A606 ,
    A607 , A608 , A609 , A610 , A611 , A612 , A613 ,
    A614 , A615 , A616 , A617 , A618 , A619 , A620 ,
    A621 , A622 , A623 , A624 , A625 , A626 , A627 ,
    A628 , A629 , A630 , A631 , A632 , A633 , A634 ,
    A635 , A636 , A637 , A638 , A639 , A640 , A641 ,
    A642 , A643 , A644 , A645 , A646 , A647 , A648 ,
    A649 , A650 , A651 , A652 , A653 , A654 , A655 ,
    A656 , A657 , A658 , A659 , A660 , A661 , A662 ,
    A663 , A664 , A665 , A666 , A667 , A668 , A669 ,
    A670 , A671 , A672 , A673 , A674 , A675 , A676 ,
    A677 , A678 , A679 , A680 , A681 , A682 , A683 ,
    A684 , A685 , A686 , A687 , A688 , A689 , A690 ,
    A691 , A692 , A693 , A694 , A695 , A696 , A697 ,
    A698 , A699 , A700 , A701 , A702 , A703 , A704 ,
    A705 , A706 , A707 , A708 , A709 , A710 , A711 ,
    A712 , A713 , A714 , A715 , A716 , A717 , A718 ,
    A719 , A720 , A721 , A722 , A723 , A724 , A725 ,
    A726 , A727 , A728 , A729 , A730 , A731 , A732 ,
    A733 , A734 , A735 , A736 , A737 , A738 , A739 ,
    A740 , A741 , A742 , A743 , A744 , A745 , A746 ,
    A747 , A748 , A749 , A750 , A751 , A752 , A753 ,
    A754 , A755 , A756 , A757 , A758 , A759 , A760 ,
    A761 , A762 , A763 , A764 , A765 , A766 , A767 ,
    A768 , A769 , A770 , A771 , A772 , A773 , A774 ,
    A775 , A776 , A777 , A778 , A779 , A780 , A781 ,
    A782 , A783 , A784 , A785 , A786 , A787 , A788 ,
    A789 , A790 , A791 , A792 , A793 , A794 , A795 ,
    A796 , A797 , A798 , A799 , A800 , A801 , A802 ,
    A803 , A804 , A805 , A806 , A807 , A808 , A809 ,
    A810 , A811 , A812 , A813 , A814 , A815 , A816 ,
    A817 , A818 , A819 , A820 , A821 , A822 , A823 ,
    A824 , A825 , A826 , A827 , A828 , A829 , A830 ,
    A831 , A832 , A833 , A834 , A835 , A836 , A837 ,
    A838 , A839 , A840 , A841 , A842 , A843 , A844 ,
    A845 , A846 , A847 , A848 , A849 , A850 , A851 ,
    A852 , A853 , A854 , A855 , A856 , A857 , A858 ,
    A859 , A860 , A861 , A862 , A863 , A864 , A865 ,
    A866 , A867 , A868 , A869 , A870 , A871 , A872 ,
    A873 , A874 , A875 , A876 , A877 , A878 , A879 ,
    A880 , A881 , A882 , A883 , A884 , A885 , A886 ,
    A887 , A888 , A889 , A890 , A891 , A892 , A893 ,
    A894 , A895 , A896 , A897 , A898 , A899 , A900 ,
    A901 , A902 , A903 , A904 , A905 , A906 , A907 ,
    A908 , A909 , A910 , A911 , A912 , A913 , A914 ,
    A915 , A916 , A917 , A918 , A919 , A920 , A921 ,
    A922 , A923 , A924 , A925 , A926 , A927 , A928 ,
    A929 , A930 , A931 , A932 , A933 , A934 , A935 ,
    A936 , A937 , A938 , A939 , A940 , A941 , A942 ,
    A943 , A944 , A945 , A946 , A947 , A948 , A949 ,
    A950 , A951 , A952 , A953 , A954 , A955 , A956 ,
    A957 , A958 , A959 , A960 , A961 , A962 , A963 ,
    A964 , A965 , A966 , A967 , A968 , A969 , A970 ,
    A971 , A972 , A973 , A974 , A975 , A976 , A977 ,
    A978 , A979 , A980 , A981 , A982 , A983 , A984 ,
    A985 , A986 , A987 , A988 , A989 , A990 , A991 ,
    A992 , A993 , A994 , A995 , A996 , A997 , A998 ,
    A999 , A1000 ;
  output maj;
  wire n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
    n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
    n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
    n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
    n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
    n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
    n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
    n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
    n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
    n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
    n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
    n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
    n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
    n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
    n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
    n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
    n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
    n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
    n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
    n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
    n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
    n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
    n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
    n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
    n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
    n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
    n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
    n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
    n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
    n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
    n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
    n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
    n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
    n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
    n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
    n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
    n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
    n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
    n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
    n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
    n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
    n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
    n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
    n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
    n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
    n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
    n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
    n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
    n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
    n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
    n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
    n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
    n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
    n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
    n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
    n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
    n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
    n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
    n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
    n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
    n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
    n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
    n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
    n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
    n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
    n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
    n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
    n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
    n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
    n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
    n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
    n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
    n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
    n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
    n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
    n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
    n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
    n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
    n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
    n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
    n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
    n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
    n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
    n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
    n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
    n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
    n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
    n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
    n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
    n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
    n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
    n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
    n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
    n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
    n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
    n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
    n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
    n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
    n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
    n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
    n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
    n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
    n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
    n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
    n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
    n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
    n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
    n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
    n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
    n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
    n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
    n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
    n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
    n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
    n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
    n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
    n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
    n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
    n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
    n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
    n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
    n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
    n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
    n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
    n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
    n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
    n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
    n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
    n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
    n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
    n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
    n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
    n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
    n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
    n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
    n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
    n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
    n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
    n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
    n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
    n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
    n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
    n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
    n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
    n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
    n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
    n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
    n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
    n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
    n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
    n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
    n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
    n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
    n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
    n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
    n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
    n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
    n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
    n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
    n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
    n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
    n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
    n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
    n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
    n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
    n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
    n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
    n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
    n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
    n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
    n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
    n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
    n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
    n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
    n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
    n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
    n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
    n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
    n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
    n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
    n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
    n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
    n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
    n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
    n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
    n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
    n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
    n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
    n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
    n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
    n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
    n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
    n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
    n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
    n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
    n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
    n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
    n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
    n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
    n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
    n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
    n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
    n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
    n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
    n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
    n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
    n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
    n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
    n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
    n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
    n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
    n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
    n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
    n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
    n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
    n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
    n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
    n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
    n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
    n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
    n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
    n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
    n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
    n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
    n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
    n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
    n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
    n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
    n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
    n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
    n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
    n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
    n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
    n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
    n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
    n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
    n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
    n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
    n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
    n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
    n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
    n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
    n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
    n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
    n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
    n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
    n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
    n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
    n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
    n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
    n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
    n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
    n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
    n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
    n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
    n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
    n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
    n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
    n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
    n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
    n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
    n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
    n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
    n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
    n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
    n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
    n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
    n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
    n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
    n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
    n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
    n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
    n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
    n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
    n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
    n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
    n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
    n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
    n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
    n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
    n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
    n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
    n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
    n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
    n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
    n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
    n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
    n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
    n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
    n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
    n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
    n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
    n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
    n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
    n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
    n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
    n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
    n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
    n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
    n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
    n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
    n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
    n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
    n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
    n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
    n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
    n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
    n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
    n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
    n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
    n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
    n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
    n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
    n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
    n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
    n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
    n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
    n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
    n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
    n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
    n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
    n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
    n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
    n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
    n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
    n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
    n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
    n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
    n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
    n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
    n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
    n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
    n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
    n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
    n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
    n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
    n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
    n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
    n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
    n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
    n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
    n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
    n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
    n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
    n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
    n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
    n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
    n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
    n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
    n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
    n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
    n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
    n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
    n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
    n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
    n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
    n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
    n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
    n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
    n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
    n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
    n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
    n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
    n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
    n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
    n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
    n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
    n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
    n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
    n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
    n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
    n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
    n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
    n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
    n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
    n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
    n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
    n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
    n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
    n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
    n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
    n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
    n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
    n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
    n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
    n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
    n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
    n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
    n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
    n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
    n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
    n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
    n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
    n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
    n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
    n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
    n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
    n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
    n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
    n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
    n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
    n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
    n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
    n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
    n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
    n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
    n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
    n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
    n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
    n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
    n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
    n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
    n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
    n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
    n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
    n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
    n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
    n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
    n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
    n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
    n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
    n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
    n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
    n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
    n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
    n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
    n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
    n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
    n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
    n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
    n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
    n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
    n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
    n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
    n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
    n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
    n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
    n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
    n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
    n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
    n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
    n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
    n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
    n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
    n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
    n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
    n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
    n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
    n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
    n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
    n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
    n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
    n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
    n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
    n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
    n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
    n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
    n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
    n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
    n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
    n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
    n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
    n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
    n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
    n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
    n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
    n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
    n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
    n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
    n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
    n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
    n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
    n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
    n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
    n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
    n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
    n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
    n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
    n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
    n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
    n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
    n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
    n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
    n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
    n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
    n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
    n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
    n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
    n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
    n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
    n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
    n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
    n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
    n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
    n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
    n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
    n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
    n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
    n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
    n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
    n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
    n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
    n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
    n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
    n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
    n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
    n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
    n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
    n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
    n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
    n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
    n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
    n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
    n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
    n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
    n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
    n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
    n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
    n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
    n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
    n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
    n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
    n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
    n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
    n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
    n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
    n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
    n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
    n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
    n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
    n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
    n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
    n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
    n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
    n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
    n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
    n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
    n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
    n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
    n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
    n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
    n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
    n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
    n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
    n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
    n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
    n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
    n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
    n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
    n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
    n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
    n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
    n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
    n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
    n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
    n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
    n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
    n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
    n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
    n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
    n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
    n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
    n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
    n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
    n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
    n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
    n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
    n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
    n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
    n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
    n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
    n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
    n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
    n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
    n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
    n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
    n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
    n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
    n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
    n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
    n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
    n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
    n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
    n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
    n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
    n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
    n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
    n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
    n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
    n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
    n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
    n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
    n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
    n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
    n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
    n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
    n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
    n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
    n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
    n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
    n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
    n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
    n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
    n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
    n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
    n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
    n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
    n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
    n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
    n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
    n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
    n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
    n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
    n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
    n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
    n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
    n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
    n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
    n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
    n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
    n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
    n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
    n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
    n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
    n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
    n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
    n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
    n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
    n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
    n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
    n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
    n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
    n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
    n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
    n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
    n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
    n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
    n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
    n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
    n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
    n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
    n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
    n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
    n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
    n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
    n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
    n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
    n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
    n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
    n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
    n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
    n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
    n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
    n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
    n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
    n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
    n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
    n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
    n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
    n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
    n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
    n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
    n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
    n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
    n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
    n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
    n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
    n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
    n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
    n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
    n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
    n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
    n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
    n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
    n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
    n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
    n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
    n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
    n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
    n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
    n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
    n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
    n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
    n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
    n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
    n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
    n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
    n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
    n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
    n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
    n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
    n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
    n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
    n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
    n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
    n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
    n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
    n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
    n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
    n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
    n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
    n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
    n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
    n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
    n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
    n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
    n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
    n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
    n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
    n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
    n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
    n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
    n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
    n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
    n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
    n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
    n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
    n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
    n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
    n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
    n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
    n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
    n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
    n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
    n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
    n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
    n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
    n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
    n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
    n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
    n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
    n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
    n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
    n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
    n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
    n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
    n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
    n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
    n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
    n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
    n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
    n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
    n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
    n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
    n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
    n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
    n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
    n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
    n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
    n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
    n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
    n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
    n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
    n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
    n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
    n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
    n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
    n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
    n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
    n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
    n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
    n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
    n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
    n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
    n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
    n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
    n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
    n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
    n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
    n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
    n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
    n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
    n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
    n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
    n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
    n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
    n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
    n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
    n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
    n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
    n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
    n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
    n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
    n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
    n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
    n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
    n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
    n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
    n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
    n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
    n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
    n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
    n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
    n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
    n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
    n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
    n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
    n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
    n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
    n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
    n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
    n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
    n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
    n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
    n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
    n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
    n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
    n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
    n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
    n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
    n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
    n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
    n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
    n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
    n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
    n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
    n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
    n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
    n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
    n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
    n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
    n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
    n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
    n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
    n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
    n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
    n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
    n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
    n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
    n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
    n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
    n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
    n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
    n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
    n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
    n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
    n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
    n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
    n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
    n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
    n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
    n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
    n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
    n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
    n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
    n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
    n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
    n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
    n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
    n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
    n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
    n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
    n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
    n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
    n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
    n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
    n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
    n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
    n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
    n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
    n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
    n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
    n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
    n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
    n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
    n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
    n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
    n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
    n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
    n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
    n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
    n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
    n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
    n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
    n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
    n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
    n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
    n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
    n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
    n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
    n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
    n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
    n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
    n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
    n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
    n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
    n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
    n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
    n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
    n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
    n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
    n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
    n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
    n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
    n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
    n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
    n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
    n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
    n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
    n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
    n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
    n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
    n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
    n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
    n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
    n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
    n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
    n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
    n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
    n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
    n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
    n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
    n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
    n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
    n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
    n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
    n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
    n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
    n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
    n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
    n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
    n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
    n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
    n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
    n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
    n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
    n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
    n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
    n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
    n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
    n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
    n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
    n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
    n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
    n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
    n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
    n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
    n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
    n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
    n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
    n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
    n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
    n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
    n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
    n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
    n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
    n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
    n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
    n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
    n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
    n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
    n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
    n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
    n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
    n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
    n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
    n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
    n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
    n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
    n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
    n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
    n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
    n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
    n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
    n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
    n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
    n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
    n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
    n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
    n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
    n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
    n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
    n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
    n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
    n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
    n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
    n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
    n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
    n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
    n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
    n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
    n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
    n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
    n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
    n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
    n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
    n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
    n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
    n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
    n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
    n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
    n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
    n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
    n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
    n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
    n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
    n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
    n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
    n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
    n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
    n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
    n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
    n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
    n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
    n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
    n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
    n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
    n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
    n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
    n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
    n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
    n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
    n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
    n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
    n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
    n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
    n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
    n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
    n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
    n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
    n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
    n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
    n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
    n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
    n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
    n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
    n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
    n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
    n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
    n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
    n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
    n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
    n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
    n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
    n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
    n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
    n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
    n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
    n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
    n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
    n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
    n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
    n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
    n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
    n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
    n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
    n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
    n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
    n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
    n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
    n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
    n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
    n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
    n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
    n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
    n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
    n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
    n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
    n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
    n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
    n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
    n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
    n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
    n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
    n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
    n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
    n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
    n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
    n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
    n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
    n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
    n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
    n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
    n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
    n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
    n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
    n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
    n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
    n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
    n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
    n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
    n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
    n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
    n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
    n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
    n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
    n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
    n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
    n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
    n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
    n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
    n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
    n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
    n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
    n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
    n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
    n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
    n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
    n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
    n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
    n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
    n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
    n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
    n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
    n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
    n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
    n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
    n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
    n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
    n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
    n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
    n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
    n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
    n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
    n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
    n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
    n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
    n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
    n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
    n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
    n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
    n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
    n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
    n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
    n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
    n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
    n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
    n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
    n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
    n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
    n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
    n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
    n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
    n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
    n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
    n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
    n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
    n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
    n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
    n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
    n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
    n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
    n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
    n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
    n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
    n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
    n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
    n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
    n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
    n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
    n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
    n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
    n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
    n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
    n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
    n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
    n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
    n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
    n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
    n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
    n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
    n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
    n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
    n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
    n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
    n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
    n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
    n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
    n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
    n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
    n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
    n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
    n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
    n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
    n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
    n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
    n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
    n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
    n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
    n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
    n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
    n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
    n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
    n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
    n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
    n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
    n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
    n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
    n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
    n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
    n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
    n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
    n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
    n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
    n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
    n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
    n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
    n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
    n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
    n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
    n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
    n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
    n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
    n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
    n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
    n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
    n14754, n14755, n14756, n14757, n14758, n14759;
  assign n1003 = A718  & A719 ;
  assign n1004 = A718  & ~A719 ;
  assign n1005 = ~A718  & A719 ;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = A720  & ~n1006;
  assign n1008 = ~n1003 & ~n1007;
  assign n1009 = A715  & A716 ;
  assign n1010 = A715  & ~A716 ;
  assign n1011 = ~A715  & A716 ;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = A717  & ~n1012;
  assign n1014 = ~n1009 & ~n1013;
  assign n1015 = n1008 & ~n1014;
  assign n1016 = ~n1008 & n1014;
  assign n1017 = A717  & ~n1010;
  assign n1018 = ~n1011 & n1017;
  assign n1019 = ~A717  & ~n1012;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = A720  & ~n1004;
  assign n1022 = ~n1005 & n1021;
  assign n1023 = ~A720  & ~n1006;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = ~n1020 & ~n1024;
  assign n1026 = ~n1016 & n1025;
  assign n1027 = ~n1015 & n1026;
  assign n1028 = ~n1015 & ~n1016;
  assign n1029 = ~n1025 & ~n1028;
  assign n1030 = ~n1027 & ~n1029;
  assign n1031 = ~n1020 & n1024;
  assign n1032 = n1020 & ~n1024;
  assign n1033 = ~n1031 & ~n1032;
  assign n1034 = n1025 & ~n1028;
  assign n1035 = ~n1008 & ~n1014;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037 = ~n1033 & ~n1036;
  assign n1038 = ~n1030 & ~n1037;
  assign n1039 = ~n1030 & ~n1036;
  assign n1040 = A724  & A725 ;
  assign n1041 = A724  & ~A725 ;
  assign n1042 = ~A724  & A725 ;
  assign n1043 = ~n1041 & ~n1042;
  assign n1044 = A726  & ~n1043;
  assign n1045 = ~n1040 & ~n1044;
  assign n1046 = A721  & A722 ;
  assign n1047 = A721  & ~A722 ;
  assign n1048 = ~A721  & A722 ;
  assign n1049 = ~n1047 & ~n1048;
  assign n1050 = A723  & ~n1049;
  assign n1051 = ~n1046 & ~n1050;
  assign n1052 = ~n1045 & n1051;
  assign n1053 = n1045 & ~n1051;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = A723  & ~n1047;
  assign n1056 = ~n1048 & n1055;
  assign n1057 = ~A723  & ~n1049;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = A726  & ~n1041;
  assign n1060 = ~n1042 & n1059;
  assign n1061 = ~A726  & ~n1043;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~n1058 & ~n1062;
  assign n1064 = ~n1054 & n1063;
  assign n1065 = ~n1045 & ~n1051;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = ~n1052 & n1063;
  assign n1068 = ~n1053 & n1067;
  assign n1069 = ~n1054 & ~n1063;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = ~n1066 & ~n1070;
  assign n1072 = ~n1058 & n1062;
  assign n1073 = n1058 & ~n1062;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = ~n1033 & ~n1074;
  assign n1076 = ~n1071 & n1075;
  assign n1077 = ~n1039 & n1076;
  assign n1078 = ~n1066 & ~n1074;
  assign n1079 = ~n1070 & ~n1078;
  assign n1080 = ~n1077 & ~n1079;
  assign n1081 = ~n1070 & n1075;
  assign n1082 = ~n1071 & n1081;
  assign n1083 = ~n1039 & ~n1078;
  assign n1084 = n1082 & n1083;
  assign n1085 = ~n1080 & ~n1084;
  assign n1086 = n1038 & ~n1085;
  assign n1087 = ~n1077 & n1079;
  assign n1088 = n1077 & ~n1079;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = ~n1038 & ~n1089;
  assign n1091 = ~n1071 & ~n1074;
  assign n1092 = ~n1033 & ~n1039;
  assign n1093 = ~n1091 & n1092;
  assign n1094 = n1091 & ~n1092;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = ~A709  & A710 ;
  assign n1097 = A709  & ~A710 ;
  assign n1098 = A711  & ~n1097;
  assign n1099 = ~n1096 & n1098;
  assign n1100 = ~n1096 & ~n1097;
  assign n1101 = ~A711  & ~n1100;
  assign n1102 = ~n1099 & ~n1101;
  assign n1103 = ~A712  & A713 ;
  assign n1104 = A712  & ~A713 ;
  assign n1105 = A714  & ~n1104;
  assign n1106 = ~n1103 & n1105;
  assign n1107 = ~n1103 & ~n1104;
  assign n1108 = ~A714  & ~n1107;
  assign n1109 = ~n1106 & ~n1108;
  assign n1110 = ~n1102 & n1109;
  assign n1111 = n1102 & ~n1109;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = A712  & A713 ;
  assign n1114 = A714  & ~n1107;
  assign n1115 = ~n1113 & ~n1114;
  assign n1116 = A709  & A710 ;
  assign n1117 = A711  & ~n1100;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = ~n1115 & n1118;
  assign n1120 = n1115 & ~n1118;
  assign n1121 = ~n1119 & ~n1120;
  assign n1122 = ~n1102 & ~n1109;
  assign n1123 = ~n1121 & n1122;
  assign n1124 = ~n1115 & ~n1118;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = ~n1119 & n1122;
  assign n1127 = ~n1120 & n1126;
  assign n1128 = ~n1121 & ~n1122;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = ~n1125 & ~n1129;
  assign n1131 = ~n1112 & ~n1130;
  assign n1132 = ~A703  & A704 ;
  assign n1133 = A703  & ~A704 ;
  assign n1134 = A705  & ~n1133;
  assign n1135 = ~n1132 & n1134;
  assign n1136 = ~n1132 & ~n1133;
  assign n1137 = ~A705  & ~n1136;
  assign n1138 = ~n1135 & ~n1137;
  assign n1139 = ~A706  & A707 ;
  assign n1140 = A706  & ~A707 ;
  assign n1141 = A708  & ~n1140;
  assign n1142 = ~n1139 & n1141;
  assign n1143 = ~n1139 & ~n1140;
  assign n1144 = ~A708  & ~n1143;
  assign n1145 = ~n1142 & ~n1144;
  assign n1146 = ~n1138 & n1145;
  assign n1147 = n1138 & ~n1145;
  assign n1148 = ~n1146 & ~n1147;
  assign n1149 = A706  & A707 ;
  assign n1150 = A708  & ~n1143;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = A703  & A704 ;
  assign n1153 = A705  & ~n1136;
  assign n1154 = ~n1152 & ~n1153;
  assign n1155 = ~n1151 & n1154;
  assign n1156 = n1151 & ~n1154;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = ~n1138 & ~n1145;
  assign n1159 = ~n1157 & n1158;
  assign n1160 = ~n1151 & ~n1154;
  assign n1161 = ~n1159 & ~n1160;
  assign n1162 = ~n1155 & n1158;
  assign n1163 = ~n1156 & n1162;
  assign n1164 = ~n1157 & ~n1158;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = ~n1161 & ~n1165;
  assign n1167 = ~n1148 & ~n1166;
  assign n1168 = ~n1131 & n1167;
  assign n1169 = n1131 & ~n1167;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = ~n1095 & ~n1170;
  assign n1172 = ~n1090 & n1171;
  assign n1173 = ~n1086 & n1172;
  assign n1174 = ~n1086 & ~n1090;
  assign n1175 = ~n1171 & ~n1174;
  assign n1176 = ~n1173 & ~n1175;
  assign n1177 = ~n1148 & ~n1161;
  assign n1178 = ~n1165 & ~n1177;
  assign n1179 = ~n1112 & ~n1148;
  assign n1180 = ~n1130 & n1179;
  assign n1181 = ~n1166 & n1180;
  assign n1182 = ~n1112 & ~n1125;
  assign n1183 = ~n1129 & ~n1182;
  assign n1184 = ~n1181 & n1183;
  assign n1185 = n1181 & ~n1183;
  assign n1186 = ~n1184 & ~n1185;
  assign n1187 = ~n1178 & ~n1186;
  assign n1188 = ~n1181 & ~n1183;
  assign n1189 = ~n1129 & n1179;
  assign n1190 = ~n1130 & n1189;
  assign n1191 = ~n1166 & ~n1182;
  assign n1192 = n1190 & n1191;
  assign n1193 = ~n1188 & ~n1192;
  assign n1194 = n1178 & ~n1193;
  assign n1195 = ~n1187 & ~n1194;
  assign n1196 = ~n1176 & n1195;
  assign n1197 = ~n1090 & ~n1171;
  assign n1198 = ~n1086 & n1197;
  assign n1199 = n1171 & ~n1174;
  assign n1200 = ~n1198 & ~n1199;
  assign n1201 = ~n1195 & ~n1200;
  assign n1202 = ~n1196 & ~n1201;
  assign n1203 = A730  & A731 ;
  assign n1204 = A730  & ~A731 ;
  assign n1205 = ~A730  & A731 ;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = A732  & ~n1206;
  assign n1208 = ~n1203 & ~n1207;
  assign n1209 = A727  & A728 ;
  assign n1210 = A727  & ~A728 ;
  assign n1211 = ~A727  & A728 ;
  assign n1212 = ~n1210 & ~n1211;
  assign n1213 = A729  & ~n1212;
  assign n1214 = ~n1209 & ~n1213;
  assign n1215 = n1208 & ~n1214;
  assign n1216 = ~n1208 & n1214;
  assign n1217 = A729  & ~n1210;
  assign n1218 = ~n1211 & n1217;
  assign n1219 = ~A729  & ~n1212;
  assign n1220 = ~n1218 & ~n1219;
  assign n1221 = A732  & ~n1204;
  assign n1222 = ~n1205 & n1221;
  assign n1223 = ~A732  & ~n1206;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = ~n1220 & ~n1224;
  assign n1226 = ~n1216 & n1225;
  assign n1227 = ~n1215 & n1226;
  assign n1228 = ~n1215 & ~n1216;
  assign n1229 = ~n1225 & ~n1228;
  assign n1230 = ~n1227 & ~n1229;
  assign n1231 = ~n1220 & n1224;
  assign n1232 = n1220 & ~n1224;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = n1225 & ~n1228;
  assign n1235 = ~n1208 & ~n1214;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = ~n1233 & ~n1236;
  assign n1238 = ~n1230 & ~n1237;
  assign n1239 = ~n1230 & ~n1236;
  assign n1240 = A736  & A737 ;
  assign n1241 = A736  & ~A737 ;
  assign n1242 = ~A736  & A737 ;
  assign n1243 = ~n1241 & ~n1242;
  assign n1244 = A738  & ~n1243;
  assign n1245 = ~n1240 & ~n1244;
  assign n1246 = A733  & A734 ;
  assign n1247 = A733  & ~A734 ;
  assign n1248 = ~A733  & A734 ;
  assign n1249 = ~n1247 & ~n1248;
  assign n1250 = A735  & ~n1249;
  assign n1251 = ~n1246 & ~n1250;
  assign n1252 = ~n1245 & n1251;
  assign n1253 = n1245 & ~n1251;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = A735  & ~n1247;
  assign n1256 = ~n1248 & n1255;
  assign n1257 = ~A735  & ~n1249;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = A738  & ~n1241;
  assign n1260 = ~n1242 & n1259;
  assign n1261 = ~A738  & ~n1243;
  assign n1262 = ~n1260 & ~n1261;
  assign n1263 = ~n1258 & ~n1262;
  assign n1264 = ~n1254 & n1263;
  assign n1265 = ~n1245 & ~n1251;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = ~n1252 & n1263;
  assign n1268 = ~n1253 & n1267;
  assign n1269 = ~n1254 & ~n1263;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = ~n1266 & ~n1270;
  assign n1272 = ~n1258 & n1262;
  assign n1273 = n1258 & ~n1262;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = ~n1233 & ~n1274;
  assign n1276 = ~n1271 & n1275;
  assign n1277 = ~n1239 & n1276;
  assign n1278 = ~n1266 & ~n1274;
  assign n1279 = ~n1270 & ~n1278;
  assign n1280 = ~n1277 & n1279;
  assign n1281 = n1277 & ~n1279;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = ~n1238 & ~n1282;
  assign n1284 = ~n1277 & ~n1279;
  assign n1285 = ~n1270 & n1275;
  assign n1286 = ~n1271 & n1285;
  assign n1287 = ~n1239 & ~n1278;
  assign n1288 = n1286 & n1287;
  assign n1289 = ~n1284 & ~n1288;
  assign n1290 = n1238 & ~n1289;
  assign n1291 = ~n1283 & ~n1290;
  assign n1292 = A742  & A743 ;
  assign n1293 = A742  & ~A743 ;
  assign n1294 = ~A742  & A743 ;
  assign n1295 = ~n1293 & ~n1294;
  assign n1296 = A744  & ~n1295;
  assign n1297 = ~n1292 & ~n1296;
  assign n1298 = A739  & A740 ;
  assign n1299 = A739  & ~A740 ;
  assign n1300 = ~A739  & A740 ;
  assign n1301 = ~n1299 & ~n1300;
  assign n1302 = A741  & ~n1301;
  assign n1303 = ~n1298 & ~n1302;
  assign n1304 = n1297 & ~n1303;
  assign n1305 = ~n1297 & n1303;
  assign n1306 = A741  & ~n1299;
  assign n1307 = ~n1300 & n1306;
  assign n1308 = ~A741  & ~n1301;
  assign n1309 = ~n1307 & ~n1308;
  assign n1310 = A744  & ~n1293;
  assign n1311 = ~n1294 & n1310;
  assign n1312 = ~A744  & ~n1295;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = ~n1309 & ~n1313;
  assign n1315 = ~n1305 & n1314;
  assign n1316 = ~n1304 & n1315;
  assign n1317 = ~n1304 & ~n1305;
  assign n1318 = ~n1314 & ~n1317;
  assign n1319 = ~n1316 & ~n1318;
  assign n1320 = ~n1309 & n1313;
  assign n1321 = n1309 & ~n1313;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = n1314 & ~n1317;
  assign n1324 = ~n1297 & ~n1303;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = ~n1322 & ~n1325;
  assign n1327 = ~n1319 & ~n1326;
  assign n1328 = ~n1319 & ~n1325;
  assign n1329 = A748  & A749 ;
  assign n1330 = A748  & ~A749 ;
  assign n1331 = ~A748  & A749 ;
  assign n1332 = ~n1330 & ~n1331;
  assign n1333 = A750  & ~n1332;
  assign n1334 = ~n1329 & ~n1333;
  assign n1335 = A745  & A746 ;
  assign n1336 = A745  & ~A746 ;
  assign n1337 = ~A745  & A746 ;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = A747  & ~n1338;
  assign n1340 = ~n1335 & ~n1339;
  assign n1341 = ~n1334 & n1340;
  assign n1342 = n1334 & ~n1340;
  assign n1343 = ~n1341 & ~n1342;
  assign n1344 = A747  & ~n1336;
  assign n1345 = ~n1337 & n1344;
  assign n1346 = ~A747  & ~n1338;
  assign n1347 = ~n1345 & ~n1346;
  assign n1348 = A750  & ~n1330;
  assign n1349 = ~n1331 & n1348;
  assign n1350 = ~A750  & ~n1332;
  assign n1351 = ~n1349 & ~n1350;
  assign n1352 = ~n1347 & ~n1351;
  assign n1353 = ~n1343 & n1352;
  assign n1354 = ~n1334 & ~n1340;
  assign n1355 = ~n1353 & ~n1354;
  assign n1356 = ~n1341 & n1352;
  assign n1357 = ~n1342 & n1356;
  assign n1358 = ~n1343 & ~n1352;
  assign n1359 = ~n1357 & ~n1358;
  assign n1360 = ~n1355 & ~n1359;
  assign n1361 = ~n1347 & n1351;
  assign n1362 = n1347 & ~n1351;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = ~n1322 & ~n1363;
  assign n1365 = ~n1360 & n1364;
  assign n1366 = ~n1328 & n1365;
  assign n1367 = ~n1355 & ~n1363;
  assign n1368 = ~n1359 & ~n1367;
  assign n1369 = ~n1366 & ~n1368;
  assign n1370 = ~n1359 & n1364;
  assign n1371 = ~n1360 & n1370;
  assign n1372 = ~n1328 & ~n1367;
  assign n1373 = n1371 & n1372;
  assign n1374 = ~n1369 & ~n1373;
  assign n1375 = n1327 & ~n1374;
  assign n1376 = ~n1366 & n1368;
  assign n1377 = n1366 & ~n1368;
  assign n1378 = ~n1376 & ~n1377;
  assign n1379 = ~n1327 & ~n1378;
  assign n1380 = ~n1360 & ~n1363;
  assign n1381 = ~n1322 & ~n1328;
  assign n1382 = ~n1380 & n1381;
  assign n1383 = n1380 & ~n1381;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = ~n1271 & ~n1274;
  assign n1386 = ~n1233 & ~n1239;
  assign n1387 = ~n1385 & n1386;
  assign n1388 = n1385 & ~n1386;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = ~n1384 & ~n1389;
  assign n1391 = ~n1379 & ~n1390;
  assign n1392 = ~n1375 & n1391;
  assign n1393 = ~n1375 & ~n1379;
  assign n1394 = n1390 & ~n1393;
  assign n1395 = ~n1392 & ~n1394;
  assign n1396 = ~n1291 & ~n1395;
  assign n1397 = ~n1379 & n1390;
  assign n1398 = ~n1375 & n1397;
  assign n1399 = ~n1390 & ~n1393;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = n1291 & ~n1400;
  assign n1402 = ~n1384 & n1389;
  assign n1403 = n1384 & ~n1389;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = ~n1095 & n1170;
  assign n1406 = n1095 & ~n1170;
  assign n1407 = ~n1405 & ~n1406;
  assign n1408 = ~n1404 & ~n1407;
  assign n1409 = ~n1401 & ~n1408;
  assign n1410 = ~n1396 & n1409;
  assign n1411 = ~n1396 & ~n1401;
  assign n1412 = n1408 & ~n1411;
  assign n1413 = ~n1410 & ~n1412;
  assign n1414 = ~n1202 & ~n1413;
  assign n1415 = ~n1401 & n1408;
  assign n1416 = ~n1396 & n1415;
  assign n1417 = ~n1408 & ~n1411;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = n1202 & ~n1418;
  assign n1420 = ~n1404 & n1407;
  assign n1421 = n1404 & ~n1407;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = ~A697  & A698 ;
  assign n1424 = A697  & ~A698 ;
  assign n1425 = A699  & ~n1424;
  assign n1426 = ~n1423 & n1425;
  assign n1427 = ~n1423 & ~n1424;
  assign n1428 = ~A699  & ~n1427;
  assign n1429 = ~n1426 & ~n1428;
  assign n1430 = ~A700  & A701 ;
  assign n1431 = A700  & ~A701 ;
  assign n1432 = A702  & ~n1431;
  assign n1433 = ~n1430 & n1432;
  assign n1434 = ~n1430 & ~n1431;
  assign n1435 = ~A702  & ~n1434;
  assign n1436 = ~n1433 & ~n1435;
  assign n1437 = ~n1429 & n1436;
  assign n1438 = n1429 & ~n1436;
  assign n1439 = ~n1437 & ~n1438;
  assign n1440 = A700  & A701 ;
  assign n1441 = A702  & ~n1434;
  assign n1442 = ~n1440 & ~n1441;
  assign n1443 = A697  & A698 ;
  assign n1444 = A699  & ~n1427;
  assign n1445 = ~n1443 & ~n1444;
  assign n1446 = ~n1442 & n1445;
  assign n1447 = n1442 & ~n1445;
  assign n1448 = ~n1446 & ~n1447;
  assign n1449 = ~n1429 & ~n1436;
  assign n1450 = ~n1448 & n1449;
  assign n1451 = ~n1442 & ~n1445;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = ~n1446 & n1449;
  assign n1454 = ~n1447 & n1453;
  assign n1455 = ~n1448 & ~n1449;
  assign n1456 = ~n1454 & ~n1455;
  assign n1457 = ~n1452 & ~n1456;
  assign n1458 = ~n1439 & ~n1457;
  assign n1459 = ~A691  & A692 ;
  assign n1460 = A691  & ~A692 ;
  assign n1461 = A693  & ~n1460;
  assign n1462 = ~n1459 & n1461;
  assign n1463 = ~n1459 & ~n1460;
  assign n1464 = ~A693  & ~n1463;
  assign n1465 = ~n1462 & ~n1464;
  assign n1466 = ~A694  & A695 ;
  assign n1467 = A694  & ~A695 ;
  assign n1468 = A696  & ~n1467;
  assign n1469 = ~n1466 & n1468;
  assign n1470 = ~n1466 & ~n1467;
  assign n1471 = ~A696  & ~n1470;
  assign n1472 = ~n1469 & ~n1471;
  assign n1473 = ~n1465 & n1472;
  assign n1474 = n1465 & ~n1472;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = A694  & A695 ;
  assign n1477 = A696  & ~n1470;
  assign n1478 = ~n1476 & ~n1477;
  assign n1479 = A691  & A692 ;
  assign n1480 = A693  & ~n1463;
  assign n1481 = ~n1479 & ~n1480;
  assign n1482 = ~n1478 & n1481;
  assign n1483 = n1478 & ~n1481;
  assign n1484 = ~n1482 & ~n1483;
  assign n1485 = ~n1465 & ~n1472;
  assign n1486 = ~n1484 & n1485;
  assign n1487 = ~n1478 & ~n1481;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = ~n1482 & n1485;
  assign n1490 = ~n1483 & n1489;
  assign n1491 = ~n1484 & ~n1485;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = ~n1488 & ~n1492;
  assign n1494 = ~n1475 & ~n1493;
  assign n1495 = ~n1458 & n1494;
  assign n1496 = n1458 & ~n1494;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = ~A685  & A686 ;
  assign n1499 = A685  & ~A686 ;
  assign n1500 = A687  & ~n1499;
  assign n1501 = ~n1498 & n1500;
  assign n1502 = ~n1498 & ~n1499;
  assign n1503 = ~A687  & ~n1502;
  assign n1504 = ~n1501 & ~n1503;
  assign n1505 = ~A688  & A689 ;
  assign n1506 = A688  & ~A689 ;
  assign n1507 = A690  & ~n1506;
  assign n1508 = ~n1505 & n1507;
  assign n1509 = ~n1505 & ~n1506;
  assign n1510 = ~A690  & ~n1509;
  assign n1511 = ~n1508 & ~n1510;
  assign n1512 = ~n1504 & n1511;
  assign n1513 = n1504 & ~n1511;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = A688  & A689 ;
  assign n1516 = A690  & ~n1509;
  assign n1517 = ~n1515 & ~n1516;
  assign n1518 = A685  & A686 ;
  assign n1519 = A687  & ~n1502;
  assign n1520 = ~n1518 & ~n1519;
  assign n1521 = ~n1517 & n1520;
  assign n1522 = n1517 & ~n1520;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = ~n1504 & ~n1511;
  assign n1525 = ~n1523 & n1524;
  assign n1526 = ~n1517 & ~n1520;
  assign n1527 = ~n1525 & ~n1526;
  assign n1528 = ~n1521 & n1524;
  assign n1529 = ~n1522 & n1528;
  assign n1530 = ~n1523 & ~n1524;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = ~n1527 & ~n1531;
  assign n1533 = ~n1514 & ~n1532;
  assign n1534 = ~A679  & A680 ;
  assign n1535 = A679  & ~A680 ;
  assign n1536 = A681  & ~n1535;
  assign n1537 = ~n1534 & n1536;
  assign n1538 = ~n1534 & ~n1535;
  assign n1539 = ~A681  & ~n1538;
  assign n1540 = ~n1537 & ~n1539;
  assign n1541 = ~A682  & A683 ;
  assign n1542 = A682  & ~A683 ;
  assign n1543 = A684  & ~n1542;
  assign n1544 = ~n1541 & n1543;
  assign n1545 = ~n1541 & ~n1542;
  assign n1546 = ~A684  & ~n1545;
  assign n1547 = ~n1544 & ~n1546;
  assign n1548 = ~n1540 & n1547;
  assign n1549 = n1540 & ~n1547;
  assign n1550 = ~n1548 & ~n1549;
  assign n1551 = A682  & A683 ;
  assign n1552 = A684  & ~n1545;
  assign n1553 = ~n1551 & ~n1552;
  assign n1554 = A679  & A680 ;
  assign n1555 = A681  & ~n1538;
  assign n1556 = ~n1554 & ~n1555;
  assign n1557 = ~n1553 & n1556;
  assign n1558 = n1553 & ~n1556;
  assign n1559 = ~n1557 & ~n1558;
  assign n1560 = ~n1540 & ~n1547;
  assign n1561 = ~n1559 & n1560;
  assign n1562 = ~n1553 & ~n1556;
  assign n1563 = ~n1561 & ~n1562;
  assign n1564 = ~n1557 & n1560;
  assign n1565 = ~n1558 & n1564;
  assign n1566 = ~n1559 & ~n1560;
  assign n1567 = ~n1565 & ~n1566;
  assign n1568 = ~n1563 & ~n1567;
  assign n1569 = ~n1550 & ~n1568;
  assign n1570 = ~n1533 & n1569;
  assign n1571 = n1533 & ~n1569;
  assign n1572 = ~n1570 & ~n1571;
  assign n1573 = ~n1497 & n1572;
  assign n1574 = n1497 & ~n1572;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = ~A673  & A674 ;
  assign n1577 = A673  & ~A674 ;
  assign n1578 = A675  & ~n1577;
  assign n1579 = ~n1576 & n1578;
  assign n1580 = ~n1576 & ~n1577;
  assign n1581 = ~A675  & ~n1580;
  assign n1582 = ~n1579 & ~n1581;
  assign n1583 = ~A676  & A677 ;
  assign n1584 = A676  & ~A677 ;
  assign n1585 = A678  & ~n1584;
  assign n1586 = ~n1583 & n1585;
  assign n1587 = ~n1583 & ~n1584;
  assign n1588 = ~A678  & ~n1587;
  assign n1589 = ~n1586 & ~n1588;
  assign n1590 = ~n1582 & n1589;
  assign n1591 = n1582 & ~n1589;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = A676  & A677 ;
  assign n1594 = A678  & ~n1587;
  assign n1595 = ~n1593 & ~n1594;
  assign n1596 = A673  & A674 ;
  assign n1597 = A675  & ~n1580;
  assign n1598 = ~n1596 & ~n1597;
  assign n1599 = ~n1595 & n1598;
  assign n1600 = n1595 & ~n1598;
  assign n1601 = ~n1599 & ~n1600;
  assign n1602 = ~n1582 & ~n1589;
  assign n1603 = ~n1601 & n1602;
  assign n1604 = ~n1595 & ~n1598;
  assign n1605 = ~n1603 & ~n1604;
  assign n1606 = ~n1599 & n1602;
  assign n1607 = ~n1600 & n1606;
  assign n1608 = ~n1601 & ~n1602;
  assign n1609 = ~n1607 & ~n1608;
  assign n1610 = ~n1605 & ~n1609;
  assign n1611 = ~n1592 & ~n1610;
  assign n1612 = ~A667  & A668 ;
  assign n1613 = A667  & ~A668 ;
  assign n1614 = A669  & ~n1613;
  assign n1615 = ~n1612 & n1614;
  assign n1616 = ~n1612 & ~n1613;
  assign n1617 = ~A669  & ~n1616;
  assign n1618 = ~n1615 & ~n1617;
  assign n1619 = ~A670  & A671 ;
  assign n1620 = A670  & ~A671 ;
  assign n1621 = A672  & ~n1620;
  assign n1622 = ~n1619 & n1621;
  assign n1623 = ~n1619 & ~n1620;
  assign n1624 = ~A672  & ~n1623;
  assign n1625 = ~n1622 & ~n1624;
  assign n1626 = ~n1618 & n1625;
  assign n1627 = n1618 & ~n1625;
  assign n1628 = ~n1626 & ~n1627;
  assign n1629 = A670  & A671 ;
  assign n1630 = A672  & ~n1623;
  assign n1631 = ~n1629 & ~n1630;
  assign n1632 = A667  & A668 ;
  assign n1633 = A669  & ~n1616;
  assign n1634 = ~n1632 & ~n1633;
  assign n1635 = ~n1631 & n1634;
  assign n1636 = n1631 & ~n1634;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = ~n1618 & ~n1625;
  assign n1639 = ~n1637 & n1638;
  assign n1640 = ~n1631 & ~n1634;
  assign n1641 = ~n1639 & ~n1640;
  assign n1642 = ~n1635 & n1638;
  assign n1643 = ~n1636 & n1642;
  assign n1644 = ~n1637 & ~n1638;
  assign n1645 = ~n1643 & ~n1644;
  assign n1646 = ~n1641 & ~n1645;
  assign n1647 = ~n1628 & ~n1646;
  assign n1648 = ~n1611 & n1647;
  assign n1649 = n1611 & ~n1647;
  assign n1650 = ~n1648 & ~n1649;
  assign n1651 = ~A661  & A662 ;
  assign n1652 = A661  & ~A662 ;
  assign n1653 = A663  & ~n1652;
  assign n1654 = ~n1651 & n1653;
  assign n1655 = ~n1651 & ~n1652;
  assign n1656 = ~A663  & ~n1655;
  assign n1657 = ~n1654 & ~n1656;
  assign n1658 = ~A664  & A665 ;
  assign n1659 = A664  & ~A665 ;
  assign n1660 = A666  & ~n1659;
  assign n1661 = ~n1658 & n1660;
  assign n1662 = ~n1658 & ~n1659;
  assign n1663 = ~A666  & ~n1662;
  assign n1664 = ~n1661 & ~n1663;
  assign n1665 = ~n1657 & n1664;
  assign n1666 = n1657 & ~n1664;
  assign n1667 = ~n1665 & ~n1666;
  assign n1668 = A664  & A665 ;
  assign n1669 = A666  & ~n1662;
  assign n1670 = ~n1668 & ~n1669;
  assign n1671 = A661  & A662 ;
  assign n1672 = A663  & ~n1655;
  assign n1673 = ~n1671 & ~n1672;
  assign n1674 = ~n1670 & n1673;
  assign n1675 = n1670 & ~n1673;
  assign n1676 = ~n1674 & ~n1675;
  assign n1677 = ~n1657 & ~n1664;
  assign n1678 = ~n1676 & n1677;
  assign n1679 = ~n1670 & ~n1673;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = ~n1674 & n1677;
  assign n1682 = ~n1675 & n1681;
  assign n1683 = ~n1676 & ~n1677;
  assign n1684 = ~n1682 & ~n1683;
  assign n1685 = ~n1680 & ~n1684;
  assign n1686 = ~n1667 & ~n1685;
  assign n1687 = ~A655  & A656 ;
  assign n1688 = A655  & ~A656 ;
  assign n1689 = A657  & ~n1688;
  assign n1690 = ~n1687 & n1689;
  assign n1691 = ~n1687 & ~n1688;
  assign n1692 = ~A657  & ~n1691;
  assign n1693 = ~n1690 & ~n1692;
  assign n1694 = ~A658  & A659 ;
  assign n1695 = A658  & ~A659 ;
  assign n1696 = A660  & ~n1695;
  assign n1697 = ~n1694 & n1696;
  assign n1698 = ~n1694 & ~n1695;
  assign n1699 = ~A660  & ~n1698;
  assign n1700 = ~n1697 & ~n1699;
  assign n1701 = ~n1693 & n1700;
  assign n1702 = n1693 & ~n1700;
  assign n1703 = ~n1701 & ~n1702;
  assign n1704 = A658  & A659 ;
  assign n1705 = A660  & ~n1698;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = A655  & A656 ;
  assign n1708 = A657  & ~n1691;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = ~n1706 & n1709;
  assign n1711 = n1706 & ~n1709;
  assign n1712 = ~n1710 & ~n1711;
  assign n1713 = ~n1693 & ~n1700;
  assign n1714 = ~n1712 & n1713;
  assign n1715 = ~n1706 & ~n1709;
  assign n1716 = ~n1714 & ~n1715;
  assign n1717 = ~n1710 & n1713;
  assign n1718 = ~n1711 & n1717;
  assign n1719 = ~n1712 & ~n1713;
  assign n1720 = ~n1718 & ~n1719;
  assign n1721 = ~n1716 & ~n1720;
  assign n1722 = ~n1703 & ~n1721;
  assign n1723 = ~n1686 & n1722;
  assign n1724 = n1686 & ~n1722;
  assign n1725 = ~n1723 & ~n1724;
  assign n1726 = ~n1650 & n1725;
  assign n1727 = n1650 & ~n1725;
  assign n1728 = ~n1726 & ~n1727;
  assign n1729 = ~n1575 & n1728;
  assign n1730 = n1575 & ~n1728;
  assign n1731 = ~n1729 & ~n1730;
  assign n1732 = ~n1422 & ~n1731;
  assign n1733 = ~n1419 & n1732;
  assign n1734 = ~n1414 & n1733;
  assign n1735 = ~n1414 & ~n1419;
  assign n1736 = ~n1732 & ~n1735;
  assign n1737 = ~n1734 & ~n1736;
  assign n1738 = ~n1550 & ~n1563;
  assign n1739 = ~n1567 & ~n1738;
  assign n1740 = ~n1514 & ~n1550;
  assign n1741 = ~n1532 & n1740;
  assign n1742 = ~n1568 & n1741;
  assign n1743 = ~n1514 & ~n1527;
  assign n1744 = ~n1531 & ~n1743;
  assign n1745 = ~n1742 & n1744;
  assign n1746 = n1742 & ~n1744;
  assign n1747 = ~n1745 & ~n1746;
  assign n1748 = ~n1739 & ~n1747;
  assign n1749 = ~n1742 & ~n1744;
  assign n1750 = ~n1531 & n1740;
  assign n1751 = ~n1532 & n1750;
  assign n1752 = ~n1568 & ~n1743;
  assign n1753 = n1751 & n1752;
  assign n1754 = ~n1749 & ~n1753;
  assign n1755 = n1739 & ~n1754;
  assign n1756 = ~n1748 & ~n1755;
  assign n1757 = ~n1475 & ~n1488;
  assign n1758 = ~n1492 & ~n1757;
  assign n1759 = ~n1439 & ~n1475;
  assign n1760 = ~n1457 & n1759;
  assign n1761 = ~n1493 & n1760;
  assign n1762 = ~n1439 & ~n1452;
  assign n1763 = ~n1456 & ~n1762;
  assign n1764 = ~n1761 & ~n1763;
  assign n1765 = ~n1456 & n1759;
  assign n1766 = ~n1457 & n1765;
  assign n1767 = ~n1493 & ~n1762;
  assign n1768 = n1766 & n1767;
  assign n1769 = ~n1764 & ~n1768;
  assign n1770 = n1758 & ~n1769;
  assign n1771 = ~n1761 & n1763;
  assign n1772 = n1761 & ~n1763;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = ~n1758 & ~n1773;
  assign n1775 = ~n1497 & ~n1572;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = ~n1770 & n1776;
  assign n1778 = ~n1770 & ~n1774;
  assign n1779 = n1775 & ~n1778;
  assign n1780 = ~n1777 & ~n1779;
  assign n1781 = ~n1756 & ~n1780;
  assign n1782 = ~n1774 & n1775;
  assign n1783 = ~n1770 & n1782;
  assign n1784 = ~n1775 & ~n1778;
  assign n1785 = ~n1783 & ~n1784;
  assign n1786 = n1756 & ~n1785;
  assign n1787 = ~n1575 & ~n1728;
  assign n1788 = ~n1786 & n1787;
  assign n1789 = ~n1781 & n1788;
  assign n1790 = ~n1781 & ~n1786;
  assign n1791 = ~n1787 & ~n1790;
  assign n1792 = ~n1789 & ~n1791;
  assign n1793 = ~n1628 & ~n1641;
  assign n1794 = ~n1645 & ~n1793;
  assign n1795 = ~n1592 & ~n1628;
  assign n1796 = ~n1610 & n1795;
  assign n1797 = ~n1646 & n1796;
  assign n1798 = ~n1592 & ~n1605;
  assign n1799 = ~n1609 & ~n1798;
  assign n1800 = ~n1797 & ~n1799;
  assign n1801 = ~n1609 & n1795;
  assign n1802 = ~n1610 & n1801;
  assign n1803 = ~n1646 & ~n1798;
  assign n1804 = n1802 & n1803;
  assign n1805 = ~n1800 & ~n1804;
  assign n1806 = n1794 & ~n1805;
  assign n1807 = ~n1797 & n1799;
  assign n1808 = n1797 & ~n1799;
  assign n1809 = ~n1807 & ~n1808;
  assign n1810 = ~n1794 & ~n1809;
  assign n1811 = ~n1650 & ~n1725;
  assign n1812 = ~n1810 & n1811;
  assign n1813 = ~n1806 & n1812;
  assign n1814 = ~n1806 & ~n1810;
  assign n1815 = ~n1811 & ~n1814;
  assign n1816 = ~n1813 & ~n1815;
  assign n1817 = ~n1703 & ~n1716;
  assign n1818 = ~n1720 & ~n1817;
  assign n1819 = ~n1667 & ~n1703;
  assign n1820 = ~n1685 & n1819;
  assign n1821 = ~n1721 & n1820;
  assign n1822 = ~n1667 & ~n1680;
  assign n1823 = ~n1684 & ~n1822;
  assign n1824 = ~n1821 & n1823;
  assign n1825 = n1821 & ~n1823;
  assign n1826 = ~n1824 & ~n1825;
  assign n1827 = ~n1818 & ~n1826;
  assign n1828 = ~n1821 & ~n1823;
  assign n1829 = ~n1684 & n1819;
  assign n1830 = ~n1685 & n1829;
  assign n1831 = ~n1721 & ~n1822;
  assign n1832 = n1830 & n1831;
  assign n1833 = ~n1828 & ~n1832;
  assign n1834 = n1818 & ~n1833;
  assign n1835 = ~n1827 & ~n1834;
  assign n1836 = ~n1816 & n1835;
  assign n1837 = ~n1810 & ~n1811;
  assign n1838 = ~n1806 & n1837;
  assign n1839 = n1811 & ~n1814;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = ~n1835 & ~n1840;
  assign n1842 = ~n1836 & ~n1841;
  assign n1843 = ~n1792 & n1842;
  assign n1844 = ~n1786 & ~n1787;
  assign n1845 = ~n1781 & n1844;
  assign n1846 = n1787 & ~n1790;
  assign n1847 = ~n1845 & ~n1846;
  assign n1848 = ~n1842 & ~n1847;
  assign n1849 = ~n1843 & ~n1848;
  assign n1850 = ~n1737 & n1849;
  assign n1851 = ~n1419 & ~n1732;
  assign n1852 = ~n1414 & n1851;
  assign n1853 = n1732 & ~n1735;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = ~n1849 & ~n1854;
  assign n1856 = ~n1850 & ~n1855;
  assign n1857 = A778  & A779 ;
  assign n1858 = A778  & ~A779 ;
  assign n1859 = ~A778  & A779 ;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = A780  & ~n1860;
  assign n1862 = ~n1857 & ~n1861;
  assign n1863 = A775  & A776 ;
  assign n1864 = A775  & ~A776 ;
  assign n1865 = ~A775  & A776 ;
  assign n1866 = ~n1864 & ~n1865;
  assign n1867 = A777  & ~n1866;
  assign n1868 = ~n1863 & ~n1867;
  assign n1869 = n1862 & ~n1868;
  assign n1870 = ~n1862 & n1868;
  assign n1871 = A777  & ~n1864;
  assign n1872 = ~n1865 & n1871;
  assign n1873 = ~A777  & ~n1866;
  assign n1874 = ~n1872 & ~n1873;
  assign n1875 = A780  & ~n1858;
  assign n1876 = ~n1859 & n1875;
  assign n1877 = ~A780  & ~n1860;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = ~n1874 & ~n1878;
  assign n1880 = ~n1870 & n1879;
  assign n1881 = ~n1869 & n1880;
  assign n1882 = ~n1869 & ~n1870;
  assign n1883 = ~n1879 & ~n1882;
  assign n1884 = ~n1881 & ~n1883;
  assign n1885 = ~n1874 & n1878;
  assign n1886 = n1874 & ~n1878;
  assign n1887 = ~n1885 & ~n1886;
  assign n1888 = n1879 & ~n1882;
  assign n1889 = ~n1862 & ~n1868;
  assign n1890 = ~n1888 & ~n1889;
  assign n1891 = ~n1887 & ~n1890;
  assign n1892 = ~n1884 & ~n1891;
  assign n1893 = ~n1884 & ~n1890;
  assign n1894 = A784  & A785 ;
  assign n1895 = A784  & ~A785 ;
  assign n1896 = ~A784  & A785 ;
  assign n1897 = ~n1895 & ~n1896;
  assign n1898 = A786  & ~n1897;
  assign n1899 = ~n1894 & ~n1898;
  assign n1900 = A781  & A782 ;
  assign n1901 = A781  & ~A782 ;
  assign n1902 = ~A781  & A782 ;
  assign n1903 = ~n1901 & ~n1902;
  assign n1904 = A783  & ~n1903;
  assign n1905 = ~n1900 & ~n1904;
  assign n1906 = ~n1899 & n1905;
  assign n1907 = n1899 & ~n1905;
  assign n1908 = ~n1906 & ~n1907;
  assign n1909 = A783  & ~n1901;
  assign n1910 = ~n1902 & n1909;
  assign n1911 = ~A783  & ~n1903;
  assign n1912 = ~n1910 & ~n1911;
  assign n1913 = A786  & ~n1895;
  assign n1914 = ~n1896 & n1913;
  assign n1915 = ~A786  & ~n1897;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = ~n1912 & ~n1916;
  assign n1918 = ~n1908 & n1917;
  assign n1919 = ~n1899 & ~n1905;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = ~n1906 & n1917;
  assign n1922 = ~n1907 & n1921;
  assign n1923 = ~n1908 & ~n1917;
  assign n1924 = ~n1922 & ~n1923;
  assign n1925 = ~n1920 & ~n1924;
  assign n1926 = ~n1912 & n1916;
  assign n1927 = n1912 & ~n1916;
  assign n1928 = ~n1926 & ~n1927;
  assign n1929 = ~n1887 & ~n1928;
  assign n1930 = ~n1925 & n1929;
  assign n1931 = ~n1893 & n1930;
  assign n1932 = ~n1920 & ~n1928;
  assign n1933 = ~n1924 & ~n1932;
  assign n1934 = ~n1931 & n1933;
  assign n1935 = n1931 & ~n1933;
  assign n1936 = ~n1934 & ~n1935;
  assign n1937 = ~n1892 & ~n1936;
  assign n1938 = ~n1931 & ~n1933;
  assign n1939 = ~n1924 & n1929;
  assign n1940 = ~n1925 & n1939;
  assign n1941 = ~n1893 & ~n1932;
  assign n1942 = n1940 & n1941;
  assign n1943 = ~n1938 & ~n1942;
  assign n1944 = n1892 & ~n1943;
  assign n1945 = ~n1937 & ~n1944;
  assign n1946 = A790  & A791 ;
  assign n1947 = A790  & ~A791 ;
  assign n1948 = ~A790  & A791 ;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = A792  & ~n1949;
  assign n1951 = ~n1946 & ~n1950;
  assign n1952 = A787  & A788 ;
  assign n1953 = A787  & ~A788 ;
  assign n1954 = ~A787  & A788 ;
  assign n1955 = ~n1953 & ~n1954;
  assign n1956 = A789  & ~n1955;
  assign n1957 = ~n1952 & ~n1956;
  assign n1958 = n1951 & ~n1957;
  assign n1959 = ~n1951 & n1957;
  assign n1960 = A789  & ~n1953;
  assign n1961 = ~n1954 & n1960;
  assign n1962 = ~A789  & ~n1955;
  assign n1963 = ~n1961 & ~n1962;
  assign n1964 = A792  & ~n1947;
  assign n1965 = ~n1948 & n1964;
  assign n1966 = ~A792  & ~n1949;
  assign n1967 = ~n1965 & ~n1966;
  assign n1968 = ~n1963 & ~n1967;
  assign n1969 = ~n1959 & n1968;
  assign n1970 = ~n1958 & n1969;
  assign n1971 = ~n1958 & ~n1959;
  assign n1972 = ~n1968 & ~n1971;
  assign n1973 = ~n1970 & ~n1972;
  assign n1974 = ~n1963 & n1967;
  assign n1975 = n1963 & ~n1967;
  assign n1976 = ~n1974 & ~n1975;
  assign n1977 = n1968 & ~n1971;
  assign n1978 = ~n1951 & ~n1957;
  assign n1979 = ~n1977 & ~n1978;
  assign n1980 = ~n1976 & ~n1979;
  assign n1981 = ~n1973 & ~n1980;
  assign n1982 = ~n1973 & ~n1979;
  assign n1983 = A796  & A797 ;
  assign n1984 = A796  & ~A797 ;
  assign n1985 = ~A796  & A797 ;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = A798  & ~n1986;
  assign n1988 = ~n1983 & ~n1987;
  assign n1989 = A793  & A794 ;
  assign n1990 = A793  & ~A794 ;
  assign n1991 = ~A793  & A794 ;
  assign n1992 = ~n1990 & ~n1991;
  assign n1993 = A795  & ~n1992;
  assign n1994 = ~n1989 & ~n1993;
  assign n1995 = ~n1988 & n1994;
  assign n1996 = n1988 & ~n1994;
  assign n1997 = ~n1995 & ~n1996;
  assign n1998 = A795  & ~n1990;
  assign n1999 = ~n1991 & n1998;
  assign n2000 = ~A795  & ~n1992;
  assign n2001 = ~n1999 & ~n2000;
  assign n2002 = A798  & ~n1984;
  assign n2003 = ~n1985 & n2002;
  assign n2004 = ~A798  & ~n1986;
  assign n2005 = ~n2003 & ~n2004;
  assign n2006 = ~n2001 & ~n2005;
  assign n2007 = ~n1997 & n2006;
  assign n2008 = ~n1988 & ~n1994;
  assign n2009 = ~n2007 & ~n2008;
  assign n2010 = ~n1995 & n2006;
  assign n2011 = ~n1996 & n2010;
  assign n2012 = ~n1997 & ~n2006;
  assign n2013 = ~n2011 & ~n2012;
  assign n2014 = ~n2009 & ~n2013;
  assign n2015 = ~n2001 & n2005;
  assign n2016 = n2001 & ~n2005;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = ~n1976 & ~n2017;
  assign n2019 = ~n2014 & n2018;
  assign n2020 = ~n1982 & n2019;
  assign n2021 = ~n2009 & ~n2017;
  assign n2022 = ~n2013 & ~n2021;
  assign n2023 = ~n2020 & ~n2022;
  assign n2024 = ~n2013 & n2018;
  assign n2025 = ~n2014 & n2024;
  assign n2026 = ~n1982 & ~n2021;
  assign n2027 = n2025 & n2026;
  assign n2028 = ~n2023 & ~n2027;
  assign n2029 = n1981 & ~n2028;
  assign n2030 = ~n2020 & n2022;
  assign n2031 = n2020 & ~n2022;
  assign n2032 = ~n2030 & ~n2031;
  assign n2033 = ~n1981 & ~n2032;
  assign n2034 = ~n2014 & ~n2017;
  assign n2035 = ~n1976 & ~n1982;
  assign n2036 = ~n2034 & n2035;
  assign n2037 = n2034 & ~n2035;
  assign n2038 = ~n2036 & ~n2037;
  assign n2039 = ~n1925 & ~n1928;
  assign n2040 = ~n1887 & ~n1893;
  assign n2041 = ~n2039 & n2040;
  assign n2042 = n2039 & ~n2040;
  assign n2043 = ~n2041 & ~n2042;
  assign n2044 = ~n2038 & ~n2043;
  assign n2045 = ~n2033 & ~n2044;
  assign n2046 = ~n2029 & n2045;
  assign n2047 = ~n2029 & ~n2033;
  assign n2048 = n2044 & ~n2047;
  assign n2049 = ~n2046 & ~n2048;
  assign n2050 = ~n1945 & ~n2049;
  assign n2051 = ~n2033 & n2044;
  assign n2052 = ~n2029 & n2051;
  assign n2053 = ~n2044 & ~n2047;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = n1945 & ~n2054;
  assign n2056 = ~n2038 & n2043;
  assign n2057 = n2038 & ~n2043;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = ~A769  & A770 ;
  assign n2060 = A769  & ~A770 ;
  assign n2061 = A771  & ~n2060;
  assign n2062 = ~n2059 & n2061;
  assign n2063 = ~n2059 & ~n2060;
  assign n2064 = ~A771  & ~n2063;
  assign n2065 = ~n2062 & ~n2064;
  assign n2066 = ~A772  & A773 ;
  assign n2067 = A772  & ~A773 ;
  assign n2068 = A774  & ~n2067;
  assign n2069 = ~n2066 & n2068;
  assign n2070 = ~n2066 & ~n2067;
  assign n2071 = ~A774  & ~n2070;
  assign n2072 = ~n2069 & ~n2071;
  assign n2073 = ~n2065 & n2072;
  assign n2074 = n2065 & ~n2072;
  assign n2075 = ~n2073 & ~n2074;
  assign n2076 = A772  & A773 ;
  assign n2077 = A774  & ~n2070;
  assign n2078 = ~n2076 & ~n2077;
  assign n2079 = A769  & A770 ;
  assign n2080 = A771  & ~n2063;
  assign n2081 = ~n2079 & ~n2080;
  assign n2082 = ~n2078 & n2081;
  assign n2083 = n2078 & ~n2081;
  assign n2084 = ~n2082 & ~n2083;
  assign n2085 = ~n2065 & ~n2072;
  assign n2086 = ~n2084 & n2085;
  assign n2087 = ~n2078 & ~n2081;
  assign n2088 = ~n2086 & ~n2087;
  assign n2089 = ~n2082 & n2085;
  assign n2090 = ~n2083 & n2089;
  assign n2091 = ~n2084 & ~n2085;
  assign n2092 = ~n2090 & ~n2091;
  assign n2093 = ~n2088 & ~n2092;
  assign n2094 = ~n2075 & ~n2093;
  assign n2095 = ~A763  & A764 ;
  assign n2096 = A763  & ~A764 ;
  assign n2097 = A765  & ~n2096;
  assign n2098 = ~n2095 & n2097;
  assign n2099 = ~n2095 & ~n2096;
  assign n2100 = ~A765  & ~n2099;
  assign n2101 = ~n2098 & ~n2100;
  assign n2102 = ~A766  & A767 ;
  assign n2103 = A766  & ~A767 ;
  assign n2104 = A768  & ~n2103;
  assign n2105 = ~n2102 & n2104;
  assign n2106 = ~n2102 & ~n2103;
  assign n2107 = ~A768  & ~n2106;
  assign n2108 = ~n2105 & ~n2107;
  assign n2109 = ~n2101 & n2108;
  assign n2110 = n2101 & ~n2108;
  assign n2111 = ~n2109 & ~n2110;
  assign n2112 = A766  & A767 ;
  assign n2113 = A768  & ~n2106;
  assign n2114 = ~n2112 & ~n2113;
  assign n2115 = A763  & A764 ;
  assign n2116 = A765  & ~n2099;
  assign n2117 = ~n2115 & ~n2116;
  assign n2118 = ~n2114 & n2117;
  assign n2119 = n2114 & ~n2117;
  assign n2120 = ~n2118 & ~n2119;
  assign n2121 = ~n2101 & ~n2108;
  assign n2122 = ~n2120 & n2121;
  assign n2123 = ~n2114 & ~n2117;
  assign n2124 = ~n2122 & ~n2123;
  assign n2125 = ~n2118 & n2121;
  assign n2126 = ~n2119 & n2125;
  assign n2127 = ~n2120 & ~n2121;
  assign n2128 = ~n2126 & ~n2127;
  assign n2129 = ~n2124 & ~n2128;
  assign n2130 = ~n2111 & ~n2129;
  assign n2131 = ~n2094 & n2130;
  assign n2132 = n2094 & ~n2130;
  assign n2133 = ~n2131 & ~n2132;
  assign n2134 = ~A757  & A758 ;
  assign n2135 = A757  & ~A758 ;
  assign n2136 = A759  & ~n2135;
  assign n2137 = ~n2134 & n2136;
  assign n2138 = ~n2134 & ~n2135;
  assign n2139 = ~A759  & ~n2138;
  assign n2140 = ~n2137 & ~n2139;
  assign n2141 = ~A760  & A761 ;
  assign n2142 = A760  & ~A761 ;
  assign n2143 = A762  & ~n2142;
  assign n2144 = ~n2141 & n2143;
  assign n2145 = ~n2141 & ~n2142;
  assign n2146 = ~A762  & ~n2145;
  assign n2147 = ~n2144 & ~n2146;
  assign n2148 = ~n2140 & n2147;
  assign n2149 = n2140 & ~n2147;
  assign n2150 = ~n2148 & ~n2149;
  assign n2151 = A760  & A761 ;
  assign n2152 = A762  & ~n2145;
  assign n2153 = ~n2151 & ~n2152;
  assign n2154 = A757  & A758 ;
  assign n2155 = A759  & ~n2138;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = ~n2153 & n2156;
  assign n2158 = n2153 & ~n2156;
  assign n2159 = ~n2157 & ~n2158;
  assign n2160 = ~n2140 & ~n2147;
  assign n2161 = ~n2159 & n2160;
  assign n2162 = ~n2153 & ~n2156;
  assign n2163 = ~n2161 & ~n2162;
  assign n2164 = ~n2157 & n2160;
  assign n2165 = ~n2158 & n2164;
  assign n2166 = ~n2159 & ~n2160;
  assign n2167 = ~n2165 & ~n2166;
  assign n2168 = ~n2163 & ~n2167;
  assign n2169 = ~n2150 & ~n2168;
  assign n2170 = ~A751  & A752 ;
  assign n2171 = A751  & ~A752 ;
  assign n2172 = A753  & ~n2171;
  assign n2173 = ~n2170 & n2172;
  assign n2174 = ~n2170 & ~n2171;
  assign n2175 = ~A753  & ~n2174;
  assign n2176 = ~n2173 & ~n2175;
  assign n2177 = ~A754  & A755 ;
  assign n2178 = A754  & ~A755 ;
  assign n2179 = A756  & ~n2178;
  assign n2180 = ~n2177 & n2179;
  assign n2181 = ~n2177 & ~n2178;
  assign n2182 = ~A756  & ~n2181;
  assign n2183 = ~n2180 & ~n2182;
  assign n2184 = ~n2176 & n2183;
  assign n2185 = n2176 & ~n2183;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = A754  & A755 ;
  assign n2188 = A756  & ~n2181;
  assign n2189 = ~n2187 & ~n2188;
  assign n2190 = A751  & A752 ;
  assign n2191 = A753  & ~n2174;
  assign n2192 = ~n2190 & ~n2191;
  assign n2193 = ~n2189 & n2192;
  assign n2194 = n2189 & ~n2192;
  assign n2195 = ~n2193 & ~n2194;
  assign n2196 = ~n2176 & ~n2183;
  assign n2197 = ~n2195 & n2196;
  assign n2198 = ~n2189 & ~n2192;
  assign n2199 = ~n2197 & ~n2198;
  assign n2200 = ~n2193 & n2196;
  assign n2201 = ~n2194 & n2200;
  assign n2202 = ~n2195 & ~n2196;
  assign n2203 = ~n2201 & ~n2202;
  assign n2204 = ~n2199 & ~n2203;
  assign n2205 = ~n2186 & ~n2204;
  assign n2206 = ~n2169 & n2205;
  assign n2207 = n2169 & ~n2205;
  assign n2208 = ~n2206 & ~n2207;
  assign n2209 = ~n2133 & n2208;
  assign n2210 = n2133 & ~n2208;
  assign n2211 = ~n2209 & ~n2210;
  assign n2212 = ~n2058 & ~n2211;
  assign n2213 = ~n2055 & n2212;
  assign n2214 = ~n2050 & n2213;
  assign n2215 = ~n2050 & ~n2055;
  assign n2216 = ~n2212 & ~n2215;
  assign n2217 = ~n2214 & ~n2216;
  assign n2218 = ~n2111 & ~n2124;
  assign n2219 = ~n2128 & ~n2218;
  assign n2220 = ~n2075 & ~n2111;
  assign n2221 = ~n2093 & n2220;
  assign n2222 = ~n2129 & n2221;
  assign n2223 = ~n2075 & ~n2088;
  assign n2224 = ~n2092 & ~n2223;
  assign n2225 = ~n2222 & ~n2224;
  assign n2226 = ~n2092 & n2220;
  assign n2227 = ~n2093 & n2226;
  assign n2228 = ~n2129 & ~n2223;
  assign n2229 = n2227 & n2228;
  assign n2230 = ~n2225 & ~n2229;
  assign n2231 = n2219 & ~n2230;
  assign n2232 = ~n2222 & n2224;
  assign n2233 = n2222 & ~n2224;
  assign n2234 = ~n2232 & ~n2233;
  assign n2235 = ~n2219 & ~n2234;
  assign n2236 = ~n2133 & ~n2208;
  assign n2237 = ~n2235 & n2236;
  assign n2238 = ~n2231 & n2237;
  assign n2239 = ~n2231 & ~n2235;
  assign n2240 = ~n2236 & ~n2239;
  assign n2241 = ~n2238 & ~n2240;
  assign n2242 = ~n2186 & ~n2199;
  assign n2243 = ~n2203 & ~n2242;
  assign n2244 = ~n2150 & ~n2186;
  assign n2245 = ~n2168 & n2244;
  assign n2246 = ~n2204 & n2245;
  assign n2247 = ~n2150 & ~n2163;
  assign n2248 = ~n2167 & ~n2247;
  assign n2249 = ~n2246 & n2248;
  assign n2250 = n2246 & ~n2248;
  assign n2251 = ~n2249 & ~n2250;
  assign n2252 = ~n2243 & ~n2251;
  assign n2253 = ~n2246 & ~n2248;
  assign n2254 = ~n2167 & n2244;
  assign n2255 = ~n2168 & n2254;
  assign n2256 = ~n2204 & ~n2247;
  assign n2257 = n2255 & n2256;
  assign n2258 = ~n2253 & ~n2257;
  assign n2259 = n2243 & ~n2258;
  assign n2260 = ~n2252 & ~n2259;
  assign n2261 = ~n2241 & n2260;
  assign n2262 = ~n2235 & ~n2236;
  assign n2263 = ~n2231 & n2262;
  assign n2264 = n2236 & ~n2239;
  assign n2265 = ~n2263 & ~n2264;
  assign n2266 = ~n2260 & ~n2265;
  assign n2267 = ~n2261 & ~n2266;
  assign n2268 = ~n2217 & n2267;
  assign n2269 = ~n2055 & ~n2212;
  assign n2270 = ~n2050 & n2269;
  assign n2271 = n2212 & ~n2215;
  assign n2272 = ~n2270 & ~n2271;
  assign n2273 = ~n2267 & ~n2272;
  assign n2274 = ~n2268 & ~n2273;
  assign n2275 = A814  & A815 ;
  assign n2276 = A814  & ~A815 ;
  assign n2277 = ~A814  & A815 ;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = A816  & ~n2278;
  assign n2280 = ~n2275 & ~n2279;
  assign n2281 = A811  & A812 ;
  assign n2282 = A811  & ~A812 ;
  assign n2283 = ~A811  & A812 ;
  assign n2284 = ~n2282 & ~n2283;
  assign n2285 = A813  & ~n2284;
  assign n2286 = ~n2281 & ~n2285;
  assign n2287 = n2280 & ~n2286;
  assign n2288 = ~n2280 & n2286;
  assign n2289 = A813  & ~n2282;
  assign n2290 = ~n2283 & n2289;
  assign n2291 = ~A813  & ~n2284;
  assign n2292 = ~n2290 & ~n2291;
  assign n2293 = A816  & ~n2276;
  assign n2294 = ~n2277 & n2293;
  assign n2295 = ~A816  & ~n2278;
  assign n2296 = ~n2294 & ~n2295;
  assign n2297 = ~n2292 & ~n2296;
  assign n2298 = ~n2288 & n2297;
  assign n2299 = ~n2287 & n2298;
  assign n2300 = ~n2287 & ~n2288;
  assign n2301 = ~n2297 & ~n2300;
  assign n2302 = ~n2299 & ~n2301;
  assign n2303 = ~n2292 & n2296;
  assign n2304 = n2292 & ~n2296;
  assign n2305 = ~n2303 & ~n2304;
  assign n2306 = n2297 & ~n2300;
  assign n2307 = ~n2280 & ~n2286;
  assign n2308 = ~n2306 & ~n2307;
  assign n2309 = ~n2305 & ~n2308;
  assign n2310 = ~n2302 & ~n2309;
  assign n2311 = ~n2302 & ~n2308;
  assign n2312 = A820  & A821 ;
  assign n2313 = A820  & ~A821 ;
  assign n2314 = ~A820  & A821 ;
  assign n2315 = ~n2313 & ~n2314;
  assign n2316 = A822  & ~n2315;
  assign n2317 = ~n2312 & ~n2316;
  assign n2318 = A817  & A818 ;
  assign n2319 = A817  & ~A818 ;
  assign n2320 = ~A817  & A818 ;
  assign n2321 = ~n2319 & ~n2320;
  assign n2322 = A819  & ~n2321;
  assign n2323 = ~n2318 & ~n2322;
  assign n2324 = ~n2317 & n2323;
  assign n2325 = n2317 & ~n2323;
  assign n2326 = ~n2324 & ~n2325;
  assign n2327 = A819  & ~n2319;
  assign n2328 = ~n2320 & n2327;
  assign n2329 = ~A819  & ~n2321;
  assign n2330 = ~n2328 & ~n2329;
  assign n2331 = A822  & ~n2313;
  assign n2332 = ~n2314 & n2331;
  assign n2333 = ~A822  & ~n2315;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = ~n2330 & ~n2334;
  assign n2336 = ~n2326 & n2335;
  assign n2337 = ~n2317 & ~n2323;
  assign n2338 = ~n2336 & ~n2337;
  assign n2339 = ~n2324 & n2335;
  assign n2340 = ~n2325 & n2339;
  assign n2341 = ~n2326 & ~n2335;
  assign n2342 = ~n2340 & ~n2341;
  assign n2343 = ~n2338 & ~n2342;
  assign n2344 = ~n2330 & n2334;
  assign n2345 = n2330 & ~n2334;
  assign n2346 = ~n2344 & ~n2345;
  assign n2347 = ~n2305 & ~n2346;
  assign n2348 = ~n2343 & n2347;
  assign n2349 = ~n2311 & n2348;
  assign n2350 = ~n2338 & ~n2346;
  assign n2351 = ~n2342 & ~n2350;
  assign n2352 = ~n2349 & ~n2351;
  assign n2353 = ~n2342 & n2347;
  assign n2354 = ~n2343 & n2353;
  assign n2355 = ~n2311 & ~n2350;
  assign n2356 = n2354 & n2355;
  assign n2357 = ~n2352 & ~n2356;
  assign n2358 = n2310 & ~n2357;
  assign n2359 = ~n2349 & n2351;
  assign n2360 = n2349 & ~n2351;
  assign n2361 = ~n2359 & ~n2360;
  assign n2362 = ~n2310 & ~n2361;
  assign n2363 = ~n2343 & ~n2346;
  assign n2364 = ~n2305 & ~n2311;
  assign n2365 = ~n2363 & n2364;
  assign n2366 = n2363 & ~n2364;
  assign n2367 = ~n2365 & ~n2366;
  assign n2368 = ~A805  & A806 ;
  assign n2369 = A805  & ~A806 ;
  assign n2370 = A807  & ~n2369;
  assign n2371 = ~n2368 & n2370;
  assign n2372 = ~n2368 & ~n2369;
  assign n2373 = ~A807  & ~n2372;
  assign n2374 = ~n2371 & ~n2373;
  assign n2375 = ~A808  & A809 ;
  assign n2376 = A808  & ~A809 ;
  assign n2377 = A810  & ~n2376;
  assign n2378 = ~n2375 & n2377;
  assign n2379 = ~n2375 & ~n2376;
  assign n2380 = ~A810  & ~n2379;
  assign n2381 = ~n2378 & ~n2380;
  assign n2382 = ~n2374 & n2381;
  assign n2383 = n2374 & ~n2381;
  assign n2384 = ~n2382 & ~n2383;
  assign n2385 = A808  & A809 ;
  assign n2386 = A810  & ~n2379;
  assign n2387 = ~n2385 & ~n2386;
  assign n2388 = A805  & A806 ;
  assign n2389 = A807  & ~n2372;
  assign n2390 = ~n2388 & ~n2389;
  assign n2391 = ~n2387 & n2390;
  assign n2392 = n2387 & ~n2390;
  assign n2393 = ~n2391 & ~n2392;
  assign n2394 = ~n2374 & ~n2381;
  assign n2395 = ~n2393 & n2394;
  assign n2396 = ~n2387 & ~n2390;
  assign n2397 = ~n2395 & ~n2396;
  assign n2398 = ~n2391 & n2394;
  assign n2399 = ~n2392 & n2398;
  assign n2400 = ~n2393 & ~n2394;
  assign n2401 = ~n2399 & ~n2400;
  assign n2402 = ~n2397 & ~n2401;
  assign n2403 = ~n2384 & ~n2402;
  assign n2404 = ~A799  & A800 ;
  assign n2405 = A799  & ~A800 ;
  assign n2406 = A801  & ~n2405;
  assign n2407 = ~n2404 & n2406;
  assign n2408 = ~n2404 & ~n2405;
  assign n2409 = ~A801  & ~n2408;
  assign n2410 = ~n2407 & ~n2409;
  assign n2411 = ~A802  & A803 ;
  assign n2412 = A802  & ~A803 ;
  assign n2413 = A804  & ~n2412;
  assign n2414 = ~n2411 & n2413;
  assign n2415 = ~n2411 & ~n2412;
  assign n2416 = ~A804  & ~n2415;
  assign n2417 = ~n2414 & ~n2416;
  assign n2418 = ~n2410 & n2417;
  assign n2419 = n2410 & ~n2417;
  assign n2420 = ~n2418 & ~n2419;
  assign n2421 = A802  & A803 ;
  assign n2422 = A804  & ~n2415;
  assign n2423 = ~n2421 & ~n2422;
  assign n2424 = A799  & A800 ;
  assign n2425 = A801  & ~n2408;
  assign n2426 = ~n2424 & ~n2425;
  assign n2427 = ~n2423 & n2426;
  assign n2428 = n2423 & ~n2426;
  assign n2429 = ~n2427 & ~n2428;
  assign n2430 = ~n2410 & ~n2417;
  assign n2431 = ~n2429 & n2430;
  assign n2432 = ~n2423 & ~n2426;
  assign n2433 = ~n2431 & ~n2432;
  assign n2434 = ~n2427 & n2430;
  assign n2435 = ~n2428 & n2434;
  assign n2436 = ~n2429 & ~n2430;
  assign n2437 = ~n2435 & ~n2436;
  assign n2438 = ~n2433 & ~n2437;
  assign n2439 = ~n2420 & ~n2438;
  assign n2440 = ~n2403 & n2439;
  assign n2441 = n2403 & ~n2439;
  assign n2442 = ~n2440 & ~n2441;
  assign n2443 = ~n2367 & ~n2442;
  assign n2444 = ~n2362 & n2443;
  assign n2445 = ~n2358 & n2444;
  assign n2446 = ~n2358 & ~n2362;
  assign n2447 = ~n2443 & ~n2446;
  assign n2448 = ~n2445 & ~n2447;
  assign n2449 = ~n2420 & ~n2433;
  assign n2450 = ~n2437 & ~n2449;
  assign n2451 = ~n2384 & ~n2420;
  assign n2452 = ~n2402 & n2451;
  assign n2453 = ~n2438 & n2452;
  assign n2454 = ~n2384 & ~n2397;
  assign n2455 = ~n2401 & ~n2454;
  assign n2456 = ~n2453 & n2455;
  assign n2457 = n2453 & ~n2455;
  assign n2458 = ~n2456 & ~n2457;
  assign n2459 = ~n2450 & ~n2458;
  assign n2460 = ~n2453 & ~n2455;
  assign n2461 = ~n2401 & n2451;
  assign n2462 = ~n2402 & n2461;
  assign n2463 = ~n2438 & ~n2454;
  assign n2464 = n2462 & n2463;
  assign n2465 = ~n2460 & ~n2464;
  assign n2466 = n2450 & ~n2465;
  assign n2467 = ~n2459 & ~n2466;
  assign n2468 = ~n2448 & n2467;
  assign n2469 = ~n2362 & ~n2443;
  assign n2470 = ~n2358 & n2469;
  assign n2471 = n2443 & ~n2446;
  assign n2472 = ~n2470 & ~n2471;
  assign n2473 = ~n2467 & ~n2472;
  assign n2474 = ~n2468 & ~n2473;
  assign n2475 = A826  & A827 ;
  assign n2476 = A826  & ~A827 ;
  assign n2477 = ~A826  & A827 ;
  assign n2478 = ~n2476 & ~n2477;
  assign n2479 = A828  & ~n2478;
  assign n2480 = ~n2475 & ~n2479;
  assign n2481 = A823  & A824 ;
  assign n2482 = A823  & ~A824 ;
  assign n2483 = ~A823  & A824 ;
  assign n2484 = ~n2482 & ~n2483;
  assign n2485 = A825  & ~n2484;
  assign n2486 = ~n2481 & ~n2485;
  assign n2487 = n2480 & ~n2486;
  assign n2488 = ~n2480 & n2486;
  assign n2489 = A825  & ~n2482;
  assign n2490 = ~n2483 & n2489;
  assign n2491 = ~A825  & ~n2484;
  assign n2492 = ~n2490 & ~n2491;
  assign n2493 = A828  & ~n2476;
  assign n2494 = ~n2477 & n2493;
  assign n2495 = ~A828  & ~n2478;
  assign n2496 = ~n2494 & ~n2495;
  assign n2497 = ~n2492 & ~n2496;
  assign n2498 = ~n2488 & n2497;
  assign n2499 = ~n2487 & n2498;
  assign n2500 = ~n2487 & ~n2488;
  assign n2501 = ~n2497 & ~n2500;
  assign n2502 = ~n2499 & ~n2501;
  assign n2503 = ~n2492 & n2496;
  assign n2504 = n2492 & ~n2496;
  assign n2505 = ~n2503 & ~n2504;
  assign n2506 = n2497 & ~n2500;
  assign n2507 = ~n2480 & ~n2486;
  assign n2508 = ~n2506 & ~n2507;
  assign n2509 = ~n2505 & ~n2508;
  assign n2510 = ~n2502 & ~n2509;
  assign n2511 = ~n2502 & ~n2508;
  assign n2512 = A832  & A833 ;
  assign n2513 = A832  & ~A833 ;
  assign n2514 = ~A832  & A833 ;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = A834  & ~n2515;
  assign n2517 = ~n2512 & ~n2516;
  assign n2518 = A829  & A830 ;
  assign n2519 = A829  & ~A830 ;
  assign n2520 = ~A829  & A830 ;
  assign n2521 = ~n2519 & ~n2520;
  assign n2522 = A831  & ~n2521;
  assign n2523 = ~n2518 & ~n2522;
  assign n2524 = ~n2517 & n2523;
  assign n2525 = n2517 & ~n2523;
  assign n2526 = ~n2524 & ~n2525;
  assign n2527 = A831  & ~n2519;
  assign n2528 = ~n2520 & n2527;
  assign n2529 = ~A831  & ~n2521;
  assign n2530 = ~n2528 & ~n2529;
  assign n2531 = A834  & ~n2513;
  assign n2532 = ~n2514 & n2531;
  assign n2533 = ~A834  & ~n2515;
  assign n2534 = ~n2532 & ~n2533;
  assign n2535 = ~n2530 & ~n2534;
  assign n2536 = ~n2526 & n2535;
  assign n2537 = ~n2517 & ~n2523;
  assign n2538 = ~n2536 & ~n2537;
  assign n2539 = ~n2524 & n2535;
  assign n2540 = ~n2525 & n2539;
  assign n2541 = ~n2526 & ~n2535;
  assign n2542 = ~n2540 & ~n2541;
  assign n2543 = ~n2538 & ~n2542;
  assign n2544 = ~n2530 & n2534;
  assign n2545 = n2530 & ~n2534;
  assign n2546 = ~n2544 & ~n2545;
  assign n2547 = ~n2505 & ~n2546;
  assign n2548 = ~n2543 & n2547;
  assign n2549 = ~n2511 & n2548;
  assign n2550 = ~n2538 & ~n2546;
  assign n2551 = ~n2542 & ~n2550;
  assign n2552 = ~n2549 & n2551;
  assign n2553 = n2549 & ~n2551;
  assign n2554 = ~n2552 & ~n2553;
  assign n2555 = ~n2510 & ~n2554;
  assign n2556 = ~n2549 & ~n2551;
  assign n2557 = ~n2542 & n2547;
  assign n2558 = ~n2543 & n2557;
  assign n2559 = ~n2511 & ~n2550;
  assign n2560 = n2558 & n2559;
  assign n2561 = ~n2556 & ~n2560;
  assign n2562 = n2510 & ~n2561;
  assign n2563 = ~n2555 & ~n2562;
  assign n2564 = A838  & A839 ;
  assign n2565 = A838  & ~A839 ;
  assign n2566 = ~A838  & A839 ;
  assign n2567 = ~n2565 & ~n2566;
  assign n2568 = A840  & ~n2567;
  assign n2569 = ~n2564 & ~n2568;
  assign n2570 = A835  & A836 ;
  assign n2571 = A835  & ~A836 ;
  assign n2572 = ~A835  & A836 ;
  assign n2573 = ~n2571 & ~n2572;
  assign n2574 = A837  & ~n2573;
  assign n2575 = ~n2570 & ~n2574;
  assign n2576 = n2569 & ~n2575;
  assign n2577 = ~n2569 & n2575;
  assign n2578 = A837  & ~n2571;
  assign n2579 = ~n2572 & n2578;
  assign n2580 = ~A837  & ~n2573;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = A840  & ~n2565;
  assign n2583 = ~n2566 & n2582;
  assign n2584 = ~A840  & ~n2567;
  assign n2585 = ~n2583 & ~n2584;
  assign n2586 = ~n2581 & ~n2585;
  assign n2587 = ~n2577 & n2586;
  assign n2588 = ~n2576 & n2587;
  assign n2589 = ~n2576 & ~n2577;
  assign n2590 = ~n2586 & ~n2589;
  assign n2591 = ~n2588 & ~n2590;
  assign n2592 = ~n2581 & n2585;
  assign n2593 = n2581 & ~n2585;
  assign n2594 = ~n2592 & ~n2593;
  assign n2595 = n2586 & ~n2589;
  assign n2596 = ~n2569 & ~n2575;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = ~n2594 & ~n2597;
  assign n2599 = ~n2591 & ~n2598;
  assign n2600 = ~n2591 & ~n2597;
  assign n2601 = A844  & A845 ;
  assign n2602 = A844  & ~A845 ;
  assign n2603 = ~A844  & A845 ;
  assign n2604 = ~n2602 & ~n2603;
  assign n2605 = A846  & ~n2604;
  assign n2606 = ~n2601 & ~n2605;
  assign n2607 = A841  & A842 ;
  assign n2608 = A841  & ~A842 ;
  assign n2609 = ~A841  & A842 ;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = A843  & ~n2610;
  assign n2612 = ~n2607 & ~n2611;
  assign n2613 = ~n2606 & n2612;
  assign n2614 = n2606 & ~n2612;
  assign n2615 = ~n2613 & ~n2614;
  assign n2616 = A843  & ~n2608;
  assign n2617 = ~n2609 & n2616;
  assign n2618 = ~A843  & ~n2610;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620 = A846  & ~n2602;
  assign n2621 = ~n2603 & n2620;
  assign n2622 = ~A846  & ~n2604;
  assign n2623 = ~n2621 & ~n2622;
  assign n2624 = ~n2619 & ~n2623;
  assign n2625 = ~n2615 & n2624;
  assign n2626 = ~n2606 & ~n2612;
  assign n2627 = ~n2625 & ~n2626;
  assign n2628 = ~n2613 & n2624;
  assign n2629 = ~n2614 & n2628;
  assign n2630 = ~n2615 & ~n2624;
  assign n2631 = ~n2629 & ~n2630;
  assign n2632 = ~n2627 & ~n2631;
  assign n2633 = ~n2619 & n2623;
  assign n2634 = n2619 & ~n2623;
  assign n2635 = ~n2633 & ~n2634;
  assign n2636 = ~n2594 & ~n2635;
  assign n2637 = ~n2632 & n2636;
  assign n2638 = ~n2600 & n2637;
  assign n2639 = ~n2627 & ~n2635;
  assign n2640 = ~n2631 & ~n2639;
  assign n2641 = ~n2638 & ~n2640;
  assign n2642 = ~n2631 & n2636;
  assign n2643 = ~n2632 & n2642;
  assign n2644 = ~n2600 & ~n2639;
  assign n2645 = n2643 & n2644;
  assign n2646 = ~n2641 & ~n2645;
  assign n2647 = n2599 & ~n2646;
  assign n2648 = ~n2638 & n2640;
  assign n2649 = n2638 & ~n2640;
  assign n2650 = ~n2648 & ~n2649;
  assign n2651 = ~n2599 & ~n2650;
  assign n2652 = ~n2632 & ~n2635;
  assign n2653 = ~n2594 & ~n2600;
  assign n2654 = ~n2652 & n2653;
  assign n2655 = n2652 & ~n2653;
  assign n2656 = ~n2654 & ~n2655;
  assign n2657 = ~n2543 & ~n2546;
  assign n2658 = ~n2505 & ~n2511;
  assign n2659 = ~n2657 & n2658;
  assign n2660 = n2657 & ~n2658;
  assign n2661 = ~n2659 & ~n2660;
  assign n2662 = ~n2656 & ~n2661;
  assign n2663 = ~n2651 & ~n2662;
  assign n2664 = ~n2647 & n2663;
  assign n2665 = ~n2647 & ~n2651;
  assign n2666 = n2662 & ~n2665;
  assign n2667 = ~n2664 & ~n2666;
  assign n2668 = ~n2563 & ~n2667;
  assign n2669 = ~n2651 & n2662;
  assign n2670 = ~n2647 & n2669;
  assign n2671 = ~n2662 & ~n2665;
  assign n2672 = ~n2670 & ~n2671;
  assign n2673 = n2563 & ~n2672;
  assign n2674 = ~n2656 & n2661;
  assign n2675 = n2656 & ~n2661;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = ~n2367 & n2442;
  assign n2678 = n2367 & ~n2442;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = ~n2676 & ~n2679;
  assign n2681 = ~n2673 & ~n2680;
  assign n2682 = ~n2668 & n2681;
  assign n2683 = ~n2668 & ~n2673;
  assign n2684 = n2680 & ~n2683;
  assign n2685 = ~n2682 & ~n2684;
  assign n2686 = ~n2474 & ~n2685;
  assign n2687 = ~n2673 & n2680;
  assign n2688 = ~n2668 & n2687;
  assign n2689 = ~n2680 & ~n2683;
  assign n2690 = ~n2688 & ~n2689;
  assign n2691 = n2474 & ~n2690;
  assign n2692 = ~n2676 & n2679;
  assign n2693 = n2676 & ~n2679;
  assign n2694 = ~n2692 & ~n2693;
  assign n2695 = ~n2058 & n2211;
  assign n2696 = n2058 & ~n2211;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = ~n2694 & ~n2697;
  assign n2699 = ~n2691 & ~n2698;
  assign n2700 = ~n2686 & n2699;
  assign n2701 = ~n2686 & ~n2691;
  assign n2702 = n2698 & ~n2701;
  assign n2703 = ~n2700 & ~n2702;
  assign n2704 = ~n2274 & ~n2703;
  assign n2705 = ~n2691 & n2698;
  assign n2706 = ~n2686 & n2705;
  assign n2707 = ~n2698 & ~n2701;
  assign n2708 = ~n2706 & ~n2707;
  assign n2709 = n2274 & ~n2708;
  assign n2710 = ~n2694 & n2697;
  assign n2711 = n2694 & ~n2697;
  assign n2712 = ~n2710 & ~n2711;
  assign n2713 = ~n1422 & n1731;
  assign n2714 = n1422 & ~n1731;
  assign n2715 = ~n2713 & ~n2714;
  assign n2716 = ~n2712 & ~n2715;
  assign n2717 = ~n2709 & ~n2716;
  assign n2718 = ~n2704 & n2717;
  assign n2719 = ~n2704 & ~n2709;
  assign n2720 = n2716 & ~n2719;
  assign n2721 = ~n2718 & ~n2720;
  assign n2722 = ~n1856 & ~n2721;
  assign n2723 = ~n2709 & n2716;
  assign n2724 = ~n2704 & n2723;
  assign n2725 = ~n2716 & ~n2719;
  assign n2726 = ~n2724 & ~n2725;
  assign n2727 = n1856 & ~n2726;
  assign n2728 = ~A469  & A470 ;
  assign n2729 = A469  & ~A470 ;
  assign n2730 = A471  & ~n2729;
  assign n2731 = ~n2728 & n2730;
  assign n2732 = ~n2728 & ~n2729;
  assign n2733 = ~A471  & ~n2732;
  assign n2734 = ~n2731 & ~n2733;
  assign n2735 = ~A472  & A473 ;
  assign n2736 = A472  & ~A473 ;
  assign n2737 = A474  & ~n2736;
  assign n2738 = ~n2735 & n2737;
  assign n2739 = ~n2735 & ~n2736;
  assign n2740 = ~A474  & ~n2739;
  assign n2741 = ~n2738 & ~n2740;
  assign n2742 = ~n2734 & n2741;
  assign n2743 = n2734 & ~n2741;
  assign n2744 = ~n2742 & ~n2743;
  assign n2745 = A472  & A473 ;
  assign n2746 = A474  & ~n2739;
  assign n2747 = ~n2745 & ~n2746;
  assign n2748 = A469  & A470 ;
  assign n2749 = A471  & ~n2732;
  assign n2750 = ~n2748 & ~n2749;
  assign n2751 = ~n2747 & n2750;
  assign n2752 = n2747 & ~n2750;
  assign n2753 = ~n2751 & ~n2752;
  assign n2754 = ~n2734 & ~n2741;
  assign n2755 = ~n2753 & n2754;
  assign n2756 = ~n2747 & ~n2750;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = ~n2751 & n2754;
  assign n2759 = ~n2752 & n2758;
  assign n2760 = ~n2753 & ~n2754;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = ~n2757 & ~n2761;
  assign n2763 = ~n2744 & ~n2762;
  assign n2764 = ~A466  & A467 ;
  assign n2765 = A466  & ~A467 ;
  assign n2766 = A468  & ~n2765;
  assign n2767 = ~n2764 & n2766;
  assign n2768 = ~n2764 & ~n2765;
  assign n2769 = ~A468  & ~n2768;
  assign n2770 = ~n2767 & ~n2769;
  assign n2771 = ~A463  & A464 ;
  assign n2772 = A463  & ~A464 ;
  assign n2773 = A465  & ~n2772;
  assign n2774 = ~n2771 & n2773;
  assign n2775 = ~n2771 & ~n2772;
  assign n2776 = ~A465  & ~n2775;
  assign n2777 = ~n2774 & ~n2776;
  assign n2778 = ~n2770 & n2777;
  assign n2779 = n2770 & ~n2777;
  assign n2780 = ~n2778 & ~n2779;
  assign n2781 = A466  & A467 ;
  assign n2782 = A468  & ~n2768;
  assign n2783 = ~n2781 & ~n2782;
  assign n2784 = A463  & A464 ;
  assign n2785 = A465  & ~n2775;
  assign n2786 = ~n2784 & ~n2785;
  assign n2787 = n2783 & ~n2786;
  assign n2788 = ~n2783 & n2786;
  assign n2789 = ~n2770 & ~n2777;
  assign n2790 = ~n2788 & n2789;
  assign n2791 = ~n2787 & n2790;
  assign n2792 = ~n2787 & ~n2788;
  assign n2793 = ~n2789 & ~n2792;
  assign n2794 = ~n2791 & ~n2793;
  assign n2795 = n2789 & ~n2792;
  assign n2796 = ~n2783 & ~n2786;
  assign n2797 = ~n2795 & ~n2796;
  assign n2798 = ~n2794 & ~n2797;
  assign n2799 = ~n2780 & ~n2798;
  assign n2800 = ~n2763 & n2799;
  assign n2801 = n2763 & ~n2799;
  assign n2802 = ~n2800 & ~n2801;
  assign n2803 = ~A481  & A482 ;
  assign n2804 = A481  & ~A482 ;
  assign n2805 = A483  & ~n2804;
  assign n2806 = ~n2803 & n2805;
  assign n2807 = ~n2803 & ~n2804;
  assign n2808 = ~A483  & ~n2807;
  assign n2809 = ~n2806 & ~n2808;
  assign n2810 = ~A484  & A485 ;
  assign n2811 = A484  & ~A485 ;
  assign n2812 = A486  & ~n2811;
  assign n2813 = ~n2810 & n2812;
  assign n2814 = ~n2810 & ~n2811;
  assign n2815 = ~A486  & ~n2814;
  assign n2816 = ~n2813 & ~n2815;
  assign n2817 = ~n2809 & n2816;
  assign n2818 = n2809 & ~n2816;
  assign n2819 = ~n2817 & ~n2818;
  assign n2820 = A484  & A485 ;
  assign n2821 = A486  & ~n2814;
  assign n2822 = ~n2820 & ~n2821;
  assign n2823 = A481  & A482 ;
  assign n2824 = A483  & ~n2807;
  assign n2825 = ~n2823 & ~n2824;
  assign n2826 = ~n2822 & n2825;
  assign n2827 = n2822 & ~n2825;
  assign n2828 = ~n2826 & ~n2827;
  assign n2829 = ~n2809 & ~n2816;
  assign n2830 = ~n2828 & n2829;
  assign n2831 = ~n2822 & ~n2825;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = ~n2826 & n2829;
  assign n2834 = ~n2827 & n2833;
  assign n2835 = ~n2828 & ~n2829;
  assign n2836 = ~n2834 & ~n2835;
  assign n2837 = ~n2832 & ~n2836;
  assign n2838 = ~n2819 & ~n2837;
  assign n2839 = ~A475  & A476 ;
  assign n2840 = A475  & ~A476 ;
  assign n2841 = A477  & ~n2840;
  assign n2842 = ~n2839 & n2841;
  assign n2843 = ~n2839 & ~n2840;
  assign n2844 = ~A477  & ~n2843;
  assign n2845 = ~n2842 & ~n2844;
  assign n2846 = ~A478  & A479 ;
  assign n2847 = A478  & ~A479 ;
  assign n2848 = A480  & ~n2847;
  assign n2849 = ~n2846 & n2848;
  assign n2850 = ~n2846 & ~n2847;
  assign n2851 = ~A480  & ~n2850;
  assign n2852 = ~n2849 & ~n2851;
  assign n2853 = ~n2845 & n2852;
  assign n2854 = n2845 & ~n2852;
  assign n2855 = ~n2853 & ~n2854;
  assign n2856 = A478  & A479 ;
  assign n2857 = A480  & ~n2850;
  assign n2858 = ~n2856 & ~n2857;
  assign n2859 = A475  & A476 ;
  assign n2860 = A477  & ~n2843;
  assign n2861 = ~n2859 & ~n2860;
  assign n2862 = ~n2858 & n2861;
  assign n2863 = n2858 & ~n2861;
  assign n2864 = ~n2862 & ~n2863;
  assign n2865 = ~n2845 & ~n2852;
  assign n2866 = ~n2864 & n2865;
  assign n2867 = ~n2858 & ~n2861;
  assign n2868 = ~n2866 & ~n2867;
  assign n2869 = ~n2862 & n2865;
  assign n2870 = ~n2863 & n2869;
  assign n2871 = ~n2864 & ~n2865;
  assign n2872 = ~n2870 & ~n2871;
  assign n2873 = ~n2868 & ~n2872;
  assign n2874 = ~n2855 & ~n2873;
  assign n2875 = ~n2838 & n2874;
  assign n2876 = n2838 & ~n2874;
  assign n2877 = ~n2875 & ~n2876;
  assign n2878 = ~n2802 & n2877;
  assign n2879 = n2802 & ~n2877;
  assign n2880 = ~n2878 & ~n2879;
  assign n2881 = ~A505  & A506 ;
  assign n2882 = A505  & ~A506 ;
  assign n2883 = A507  & ~n2882;
  assign n2884 = ~n2881 & n2883;
  assign n2885 = ~n2881 & ~n2882;
  assign n2886 = ~A507  & ~n2885;
  assign n2887 = ~n2884 & ~n2886;
  assign n2888 = ~A508  & A509 ;
  assign n2889 = A508  & ~A509 ;
  assign n2890 = A510  & ~n2889;
  assign n2891 = ~n2888 & n2890;
  assign n2892 = ~n2888 & ~n2889;
  assign n2893 = ~A510  & ~n2892;
  assign n2894 = ~n2891 & ~n2893;
  assign n2895 = ~n2887 & n2894;
  assign n2896 = n2887 & ~n2894;
  assign n2897 = ~n2895 & ~n2896;
  assign n2898 = A508  & A509 ;
  assign n2899 = A510  & ~n2892;
  assign n2900 = ~n2898 & ~n2899;
  assign n2901 = A505  & A506 ;
  assign n2902 = A507  & ~n2885;
  assign n2903 = ~n2901 & ~n2902;
  assign n2904 = ~n2900 & n2903;
  assign n2905 = n2900 & ~n2903;
  assign n2906 = ~n2904 & ~n2905;
  assign n2907 = ~n2887 & ~n2894;
  assign n2908 = ~n2906 & n2907;
  assign n2909 = ~n2900 & ~n2903;
  assign n2910 = ~n2908 & ~n2909;
  assign n2911 = ~n2904 & n2907;
  assign n2912 = ~n2905 & n2911;
  assign n2913 = ~n2906 & ~n2907;
  assign n2914 = ~n2912 & ~n2913;
  assign n2915 = ~n2910 & ~n2914;
  assign n2916 = ~n2897 & ~n2915;
  assign n2917 = ~A499  & A500 ;
  assign n2918 = A499  & ~A500 ;
  assign n2919 = A501  & ~n2918;
  assign n2920 = ~n2917 & n2919;
  assign n2921 = ~n2917 & ~n2918;
  assign n2922 = ~A501  & ~n2921;
  assign n2923 = ~n2920 & ~n2922;
  assign n2924 = ~A502  & A503 ;
  assign n2925 = A502  & ~A503 ;
  assign n2926 = A504  & ~n2925;
  assign n2927 = ~n2924 & n2926;
  assign n2928 = ~n2924 & ~n2925;
  assign n2929 = ~A504  & ~n2928;
  assign n2930 = ~n2927 & ~n2929;
  assign n2931 = ~n2923 & n2930;
  assign n2932 = n2923 & ~n2930;
  assign n2933 = ~n2931 & ~n2932;
  assign n2934 = A502  & A503 ;
  assign n2935 = A504  & ~n2928;
  assign n2936 = ~n2934 & ~n2935;
  assign n2937 = A499  & A500 ;
  assign n2938 = A501  & ~n2921;
  assign n2939 = ~n2937 & ~n2938;
  assign n2940 = ~n2936 & n2939;
  assign n2941 = n2936 & ~n2939;
  assign n2942 = ~n2940 & ~n2941;
  assign n2943 = ~n2923 & ~n2930;
  assign n2944 = ~n2942 & n2943;
  assign n2945 = ~n2936 & ~n2939;
  assign n2946 = ~n2944 & ~n2945;
  assign n2947 = ~n2940 & n2943;
  assign n2948 = ~n2941 & n2947;
  assign n2949 = ~n2942 & ~n2943;
  assign n2950 = ~n2948 & ~n2949;
  assign n2951 = ~n2946 & ~n2950;
  assign n2952 = ~n2933 & ~n2951;
  assign n2953 = ~n2916 & n2952;
  assign n2954 = n2916 & ~n2952;
  assign n2955 = ~n2953 & ~n2954;
  assign n2956 = ~A493  & A494 ;
  assign n2957 = A493  & ~A494 ;
  assign n2958 = A495  & ~n2957;
  assign n2959 = ~n2956 & n2958;
  assign n2960 = ~n2956 & ~n2957;
  assign n2961 = ~A495  & ~n2960;
  assign n2962 = ~n2959 & ~n2961;
  assign n2963 = ~A496  & A497 ;
  assign n2964 = A496  & ~A497 ;
  assign n2965 = A498  & ~n2964;
  assign n2966 = ~n2963 & n2965;
  assign n2967 = ~n2963 & ~n2964;
  assign n2968 = ~A498  & ~n2967;
  assign n2969 = ~n2966 & ~n2968;
  assign n2970 = ~n2962 & n2969;
  assign n2971 = n2962 & ~n2969;
  assign n2972 = ~n2970 & ~n2971;
  assign n2973 = A496  & A497 ;
  assign n2974 = A498  & ~n2967;
  assign n2975 = ~n2973 & ~n2974;
  assign n2976 = A493  & A494 ;
  assign n2977 = A495  & ~n2960;
  assign n2978 = ~n2976 & ~n2977;
  assign n2979 = ~n2975 & n2978;
  assign n2980 = n2975 & ~n2978;
  assign n2981 = ~n2979 & ~n2980;
  assign n2982 = ~n2962 & ~n2969;
  assign n2983 = ~n2981 & n2982;
  assign n2984 = ~n2975 & ~n2978;
  assign n2985 = ~n2983 & ~n2984;
  assign n2986 = ~n2979 & n2982;
  assign n2987 = ~n2980 & n2986;
  assign n2988 = ~n2981 & ~n2982;
  assign n2989 = ~n2987 & ~n2988;
  assign n2990 = ~n2985 & ~n2989;
  assign n2991 = ~n2972 & ~n2990;
  assign n2992 = ~A487  & A488 ;
  assign n2993 = A487  & ~A488 ;
  assign n2994 = A489  & ~n2993;
  assign n2995 = ~n2992 & n2994;
  assign n2996 = ~n2992 & ~n2993;
  assign n2997 = ~A489  & ~n2996;
  assign n2998 = ~n2995 & ~n2997;
  assign n2999 = ~A490  & A491 ;
  assign n3000 = A490  & ~A491 ;
  assign n3001 = A492  & ~n3000;
  assign n3002 = ~n2999 & n3001;
  assign n3003 = ~n2999 & ~n3000;
  assign n3004 = ~A492  & ~n3003;
  assign n3005 = ~n3002 & ~n3004;
  assign n3006 = ~n2998 & n3005;
  assign n3007 = n2998 & ~n3005;
  assign n3008 = ~n3006 & ~n3007;
  assign n3009 = A490  & A491 ;
  assign n3010 = A492  & ~n3003;
  assign n3011 = ~n3009 & ~n3010;
  assign n3012 = A487  & A488 ;
  assign n3013 = A489  & ~n2996;
  assign n3014 = ~n3012 & ~n3013;
  assign n3015 = ~n3011 & n3014;
  assign n3016 = n3011 & ~n3014;
  assign n3017 = ~n3015 & ~n3016;
  assign n3018 = ~n2998 & ~n3005;
  assign n3019 = ~n3017 & n3018;
  assign n3020 = ~n3011 & ~n3014;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = ~n3015 & n3018;
  assign n3023 = ~n3016 & n3022;
  assign n3024 = ~n3017 & ~n3018;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = ~n3021 & ~n3025;
  assign n3027 = ~n3008 & ~n3026;
  assign n3028 = ~n2991 & n3027;
  assign n3029 = n2991 & ~n3027;
  assign n3030 = ~n3028 & ~n3029;
  assign n3031 = ~n2955 & n3030;
  assign n3032 = n2955 & ~n3030;
  assign n3033 = ~n3031 & ~n3032;
  assign n3034 = ~n2880 & n3033;
  assign n3035 = n2880 & ~n3033;
  assign n3036 = ~n3034 & ~n3035;
  assign n3037 = ~A553  & A554 ;
  assign n3038 = A553  & ~A554 ;
  assign n3039 = A555  & ~n3038;
  assign n3040 = ~n3037 & n3039;
  assign n3041 = ~n3037 & ~n3038;
  assign n3042 = ~A555  & ~n3041;
  assign n3043 = ~n3040 & ~n3042;
  assign n3044 = ~A556  & A557 ;
  assign n3045 = A556  & ~A557 ;
  assign n3046 = A558  & ~n3045;
  assign n3047 = ~n3044 & n3046;
  assign n3048 = ~n3044 & ~n3045;
  assign n3049 = ~A558  & ~n3048;
  assign n3050 = ~n3047 & ~n3049;
  assign n3051 = ~n3043 & n3050;
  assign n3052 = n3043 & ~n3050;
  assign n3053 = ~n3051 & ~n3052;
  assign n3054 = A556  & A557 ;
  assign n3055 = A558  & ~n3048;
  assign n3056 = ~n3054 & ~n3055;
  assign n3057 = A553  & A554 ;
  assign n3058 = A555  & ~n3041;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = ~n3056 & n3059;
  assign n3061 = n3056 & ~n3059;
  assign n3062 = ~n3060 & ~n3061;
  assign n3063 = ~n3043 & ~n3050;
  assign n3064 = ~n3062 & n3063;
  assign n3065 = ~n3056 & ~n3059;
  assign n3066 = ~n3064 & ~n3065;
  assign n3067 = ~n3060 & n3063;
  assign n3068 = ~n3061 & n3067;
  assign n3069 = ~n3062 & ~n3063;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = ~n3066 & ~n3070;
  assign n3072 = ~n3053 & ~n3071;
  assign n3073 = ~A547  & A548 ;
  assign n3074 = A547  & ~A548 ;
  assign n3075 = A549  & ~n3074;
  assign n3076 = ~n3073 & n3075;
  assign n3077 = ~n3073 & ~n3074;
  assign n3078 = ~A549  & ~n3077;
  assign n3079 = ~n3076 & ~n3078;
  assign n3080 = ~A550  & A551 ;
  assign n3081 = A550  & ~A551 ;
  assign n3082 = A552  & ~n3081;
  assign n3083 = ~n3080 & n3082;
  assign n3084 = ~n3080 & ~n3081;
  assign n3085 = ~A552  & ~n3084;
  assign n3086 = ~n3083 & ~n3085;
  assign n3087 = ~n3079 & n3086;
  assign n3088 = n3079 & ~n3086;
  assign n3089 = ~n3087 & ~n3088;
  assign n3090 = A550  & A551 ;
  assign n3091 = A552  & ~n3084;
  assign n3092 = ~n3090 & ~n3091;
  assign n3093 = A547  & A548 ;
  assign n3094 = A549  & ~n3077;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = ~n3092 & n3095;
  assign n3097 = n3092 & ~n3095;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = ~n3079 & ~n3086;
  assign n3100 = ~n3098 & n3099;
  assign n3101 = ~n3092 & ~n3095;
  assign n3102 = ~n3100 & ~n3101;
  assign n3103 = ~n3096 & n3099;
  assign n3104 = ~n3097 & n3103;
  assign n3105 = ~n3098 & ~n3099;
  assign n3106 = ~n3104 & ~n3105;
  assign n3107 = ~n3102 & ~n3106;
  assign n3108 = ~n3089 & ~n3107;
  assign n3109 = ~n3072 & n3108;
  assign n3110 = n3072 & ~n3108;
  assign n3111 = ~n3109 & ~n3110;
  assign n3112 = ~A541  & A542 ;
  assign n3113 = A541  & ~A542 ;
  assign n3114 = A543  & ~n3113;
  assign n3115 = ~n3112 & n3114;
  assign n3116 = ~n3112 & ~n3113;
  assign n3117 = ~A543  & ~n3116;
  assign n3118 = ~n3115 & ~n3117;
  assign n3119 = ~A544  & A545 ;
  assign n3120 = A544  & ~A545 ;
  assign n3121 = A546  & ~n3120;
  assign n3122 = ~n3119 & n3121;
  assign n3123 = ~n3119 & ~n3120;
  assign n3124 = ~A546  & ~n3123;
  assign n3125 = ~n3122 & ~n3124;
  assign n3126 = ~n3118 & n3125;
  assign n3127 = n3118 & ~n3125;
  assign n3128 = ~n3126 & ~n3127;
  assign n3129 = A544  & A545 ;
  assign n3130 = A546  & ~n3123;
  assign n3131 = ~n3129 & ~n3130;
  assign n3132 = A541  & A542 ;
  assign n3133 = A543  & ~n3116;
  assign n3134 = ~n3132 & ~n3133;
  assign n3135 = ~n3131 & n3134;
  assign n3136 = n3131 & ~n3134;
  assign n3137 = ~n3135 & ~n3136;
  assign n3138 = ~n3118 & ~n3125;
  assign n3139 = ~n3137 & n3138;
  assign n3140 = ~n3131 & ~n3134;
  assign n3141 = ~n3139 & ~n3140;
  assign n3142 = ~n3135 & n3138;
  assign n3143 = ~n3136 & n3142;
  assign n3144 = ~n3137 & ~n3138;
  assign n3145 = ~n3143 & ~n3144;
  assign n3146 = ~n3141 & ~n3145;
  assign n3147 = ~n3128 & ~n3146;
  assign n3148 = ~A535  & A536 ;
  assign n3149 = A535  & ~A536 ;
  assign n3150 = A537  & ~n3149;
  assign n3151 = ~n3148 & n3150;
  assign n3152 = ~n3148 & ~n3149;
  assign n3153 = ~A537  & ~n3152;
  assign n3154 = ~n3151 & ~n3153;
  assign n3155 = ~A538  & A539 ;
  assign n3156 = A538  & ~A539 ;
  assign n3157 = A540  & ~n3156;
  assign n3158 = ~n3155 & n3157;
  assign n3159 = ~n3155 & ~n3156;
  assign n3160 = ~A540  & ~n3159;
  assign n3161 = ~n3158 & ~n3160;
  assign n3162 = ~n3154 & n3161;
  assign n3163 = n3154 & ~n3161;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = A538  & A539 ;
  assign n3166 = A540  & ~n3159;
  assign n3167 = ~n3165 & ~n3166;
  assign n3168 = A535  & A536 ;
  assign n3169 = A537  & ~n3152;
  assign n3170 = ~n3168 & ~n3169;
  assign n3171 = ~n3167 & n3170;
  assign n3172 = n3167 & ~n3170;
  assign n3173 = ~n3171 & ~n3172;
  assign n3174 = ~n3154 & ~n3161;
  assign n3175 = ~n3173 & n3174;
  assign n3176 = ~n3167 & ~n3170;
  assign n3177 = ~n3175 & ~n3176;
  assign n3178 = ~n3171 & n3174;
  assign n3179 = ~n3172 & n3178;
  assign n3180 = ~n3173 & ~n3174;
  assign n3181 = ~n3179 & ~n3180;
  assign n3182 = ~n3177 & ~n3181;
  assign n3183 = ~n3164 & ~n3182;
  assign n3184 = ~n3147 & n3183;
  assign n3185 = n3147 & ~n3183;
  assign n3186 = ~n3184 & ~n3185;
  assign n3187 = ~n3111 & n3186;
  assign n3188 = n3111 & ~n3186;
  assign n3189 = ~n3187 & ~n3188;
  assign n3190 = ~A529  & A530 ;
  assign n3191 = A529  & ~A530 ;
  assign n3192 = A531  & ~n3191;
  assign n3193 = ~n3190 & n3192;
  assign n3194 = ~n3190 & ~n3191;
  assign n3195 = ~A531  & ~n3194;
  assign n3196 = ~n3193 & ~n3195;
  assign n3197 = ~A532  & A533 ;
  assign n3198 = A532  & ~A533 ;
  assign n3199 = A534  & ~n3198;
  assign n3200 = ~n3197 & n3199;
  assign n3201 = ~n3197 & ~n3198;
  assign n3202 = ~A534  & ~n3201;
  assign n3203 = ~n3200 & ~n3202;
  assign n3204 = ~n3196 & n3203;
  assign n3205 = n3196 & ~n3203;
  assign n3206 = ~n3204 & ~n3205;
  assign n3207 = A532  & A533 ;
  assign n3208 = A534  & ~n3201;
  assign n3209 = ~n3207 & ~n3208;
  assign n3210 = A529  & A530 ;
  assign n3211 = A531  & ~n3194;
  assign n3212 = ~n3210 & ~n3211;
  assign n3213 = ~n3209 & n3212;
  assign n3214 = n3209 & ~n3212;
  assign n3215 = ~n3213 & ~n3214;
  assign n3216 = ~n3196 & ~n3203;
  assign n3217 = ~n3215 & n3216;
  assign n3218 = ~n3209 & ~n3212;
  assign n3219 = ~n3217 & ~n3218;
  assign n3220 = ~n3213 & n3216;
  assign n3221 = ~n3214 & n3220;
  assign n3222 = ~n3215 & ~n3216;
  assign n3223 = ~n3221 & ~n3222;
  assign n3224 = ~n3219 & ~n3223;
  assign n3225 = ~n3206 & ~n3224;
  assign n3226 = ~A523  & A524 ;
  assign n3227 = A523  & ~A524 ;
  assign n3228 = A525  & ~n3227;
  assign n3229 = ~n3226 & n3228;
  assign n3230 = ~n3226 & ~n3227;
  assign n3231 = ~A525  & ~n3230;
  assign n3232 = ~n3229 & ~n3231;
  assign n3233 = ~A526  & A527 ;
  assign n3234 = A526  & ~A527 ;
  assign n3235 = A528  & ~n3234;
  assign n3236 = ~n3233 & n3235;
  assign n3237 = ~n3233 & ~n3234;
  assign n3238 = ~A528  & ~n3237;
  assign n3239 = ~n3236 & ~n3238;
  assign n3240 = ~n3232 & n3239;
  assign n3241 = n3232 & ~n3239;
  assign n3242 = ~n3240 & ~n3241;
  assign n3243 = A526  & A527 ;
  assign n3244 = A528  & ~n3237;
  assign n3245 = ~n3243 & ~n3244;
  assign n3246 = A523  & A524 ;
  assign n3247 = A525  & ~n3230;
  assign n3248 = ~n3246 & ~n3247;
  assign n3249 = ~n3245 & n3248;
  assign n3250 = n3245 & ~n3248;
  assign n3251 = ~n3249 & ~n3250;
  assign n3252 = ~n3232 & ~n3239;
  assign n3253 = ~n3251 & n3252;
  assign n3254 = ~n3245 & ~n3248;
  assign n3255 = ~n3253 & ~n3254;
  assign n3256 = ~n3249 & n3252;
  assign n3257 = ~n3250 & n3256;
  assign n3258 = ~n3251 & ~n3252;
  assign n3259 = ~n3257 & ~n3258;
  assign n3260 = ~n3255 & ~n3259;
  assign n3261 = ~n3242 & ~n3260;
  assign n3262 = ~n3225 & n3261;
  assign n3263 = n3225 & ~n3261;
  assign n3264 = ~n3262 & ~n3263;
  assign n3265 = ~A517  & A518 ;
  assign n3266 = A517  & ~A518 ;
  assign n3267 = A519  & ~n3266;
  assign n3268 = ~n3265 & n3267;
  assign n3269 = ~n3265 & ~n3266;
  assign n3270 = ~A519  & ~n3269;
  assign n3271 = ~n3268 & ~n3270;
  assign n3272 = ~A520  & A521 ;
  assign n3273 = A520  & ~A521 ;
  assign n3274 = A522  & ~n3273;
  assign n3275 = ~n3272 & n3274;
  assign n3276 = ~n3272 & ~n3273;
  assign n3277 = ~A522  & ~n3276;
  assign n3278 = ~n3275 & ~n3277;
  assign n3279 = ~n3271 & n3278;
  assign n3280 = n3271 & ~n3278;
  assign n3281 = ~n3279 & ~n3280;
  assign n3282 = A520  & A521 ;
  assign n3283 = A522  & ~n3276;
  assign n3284 = ~n3282 & ~n3283;
  assign n3285 = A517  & A518 ;
  assign n3286 = A519  & ~n3269;
  assign n3287 = ~n3285 & ~n3286;
  assign n3288 = ~n3284 & n3287;
  assign n3289 = n3284 & ~n3287;
  assign n3290 = ~n3288 & ~n3289;
  assign n3291 = ~n3271 & ~n3278;
  assign n3292 = ~n3290 & n3291;
  assign n3293 = ~n3284 & ~n3287;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = ~n3288 & n3291;
  assign n3296 = ~n3289 & n3295;
  assign n3297 = ~n3290 & ~n3291;
  assign n3298 = ~n3296 & ~n3297;
  assign n3299 = ~n3294 & ~n3298;
  assign n3300 = ~n3281 & ~n3299;
  assign n3301 = ~A511  & A512 ;
  assign n3302 = A511  & ~A512 ;
  assign n3303 = A513  & ~n3302;
  assign n3304 = ~n3301 & n3303;
  assign n3305 = ~n3301 & ~n3302;
  assign n3306 = ~A513  & ~n3305;
  assign n3307 = ~n3304 & ~n3306;
  assign n3308 = ~A514  & A515 ;
  assign n3309 = A514  & ~A515 ;
  assign n3310 = A516  & ~n3309;
  assign n3311 = ~n3308 & n3310;
  assign n3312 = ~n3308 & ~n3309;
  assign n3313 = ~A516  & ~n3312;
  assign n3314 = ~n3311 & ~n3313;
  assign n3315 = ~n3307 & n3314;
  assign n3316 = n3307 & ~n3314;
  assign n3317 = ~n3315 & ~n3316;
  assign n3318 = A514  & A515 ;
  assign n3319 = A516  & ~n3312;
  assign n3320 = ~n3318 & ~n3319;
  assign n3321 = A511  & A512 ;
  assign n3322 = A513  & ~n3305;
  assign n3323 = ~n3321 & ~n3322;
  assign n3324 = ~n3320 & n3323;
  assign n3325 = n3320 & ~n3323;
  assign n3326 = ~n3324 & ~n3325;
  assign n3327 = ~n3307 & ~n3314;
  assign n3328 = ~n3326 & n3327;
  assign n3329 = ~n3320 & ~n3323;
  assign n3330 = ~n3328 & ~n3329;
  assign n3331 = ~n3324 & n3327;
  assign n3332 = ~n3325 & n3331;
  assign n3333 = ~n3326 & ~n3327;
  assign n3334 = ~n3332 & ~n3333;
  assign n3335 = ~n3330 & ~n3334;
  assign n3336 = ~n3317 & ~n3335;
  assign n3337 = ~n3300 & n3336;
  assign n3338 = n3300 & ~n3336;
  assign n3339 = ~n3337 & ~n3338;
  assign n3340 = ~n3264 & n3339;
  assign n3341 = n3264 & ~n3339;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = ~n3189 & n3342;
  assign n3344 = n3189 & ~n3342;
  assign n3345 = ~n3343 & ~n3344;
  assign n3346 = ~n3036 & n3345;
  assign n3347 = n3036 & ~n3345;
  assign n3348 = ~n3346 & ~n3347;
  assign n3349 = ~A649  & A650 ;
  assign n3350 = A649  & ~A650 ;
  assign n3351 = A651  & ~n3350;
  assign n3352 = ~n3349 & n3351;
  assign n3353 = ~n3349 & ~n3350;
  assign n3354 = ~A651  & ~n3353;
  assign n3355 = ~n3352 & ~n3354;
  assign n3356 = ~A652  & A653 ;
  assign n3357 = A652  & ~A653 ;
  assign n3358 = A654  & ~n3357;
  assign n3359 = ~n3356 & n3358;
  assign n3360 = ~n3356 & ~n3357;
  assign n3361 = ~A654  & ~n3360;
  assign n3362 = ~n3359 & ~n3361;
  assign n3363 = ~n3355 & n3362;
  assign n3364 = n3355 & ~n3362;
  assign n3365 = ~n3363 & ~n3364;
  assign n3366 = A652  & A653 ;
  assign n3367 = A654  & ~n3360;
  assign n3368 = ~n3366 & ~n3367;
  assign n3369 = A649  & A650 ;
  assign n3370 = A651  & ~n3353;
  assign n3371 = ~n3369 & ~n3370;
  assign n3372 = ~n3368 & n3371;
  assign n3373 = n3368 & ~n3371;
  assign n3374 = ~n3372 & ~n3373;
  assign n3375 = ~n3355 & ~n3362;
  assign n3376 = ~n3374 & n3375;
  assign n3377 = ~n3368 & ~n3371;
  assign n3378 = ~n3376 & ~n3377;
  assign n3379 = ~n3372 & n3375;
  assign n3380 = ~n3373 & n3379;
  assign n3381 = ~n3374 & ~n3375;
  assign n3382 = ~n3380 & ~n3381;
  assign n3383 = ~n3378 & ~n3382;
  assign n3384 = ~n3365 & ~n3383;
  assign n3385 = ~A643  & A644 ;
  assign n3386 = A643  & ~A644 ;
  assign n3387 = A645  & ~n3386;
  assign n3388 = ~n3385 & n3387;
  assign n3389 = ~n3385 & ~n3386;
  assign n3390 = ~A645  & ~n3389;
  assign n3391 = ~n3388 & ~n3390;
  assign n3392 = ~A646  & A647 ;
  assign n3393 = A646  & ~A647 ;
  assign n3394 = A648  & ~n3393;
  assign n3395 = ~n3392 & n3394;
  assign n3396 = ~n3392 & ~n3393;
  assign n3397 = ~A648  & ~n3396;
  assign n3398 = ~n3395 & ~n3397;
  assign n3399 = ~n3391 & n3398;
  assign n3400 = n3391 & ~n3398;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = A646  & A647 ;
  assign n3403 = A648  & ~n3396;
  assign n3404 = ~n3402 & ~n3403;
  assign n3405 = A643  & A644 ;
  assign n3406 = A645  & ~n3389;
  assign n3407 = ~n3405 & ~n3406;
  assign n3408 = ~n3404 & n3407;
  assign n3409 = n3404 & ~n3407;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = ~n3391 & ~n3398;
  assign n3412 = ~n3410 & n3411;
  assign n3413 = ~n3404 & ~n3407;
  assign n3414 = ~n3412 & ~n3413;
  assign n3415 = ~n3408 & n3411;
  assign n3416 = ~n3409 & n3415;
  assign n3417 = ~n3410 & ~n3411;
  assign n3418 = ~n3416 & ~n3417;
  assign n3419 = ~n3414 & ~n3418;
  assign n3420 = ~n3401 & ~n3419;
  assign n3421 = ~n3384 & n3420;
  assign n3422 = n3384 & ~n3420;
  assign n3423 = ~n3421 & ~n3422;
  assign n3424 = ~A637  & A638 ;
  assign n3425 = A637  & ~A638 ;
  assign n3426 = A639  & ~n3425;
  assign n3427 = ~n3424 & n3426;
  assign n3428 = ~n3424 & ~n3425;
  assign n3429 = ~A639  & ~n3428;
  assign n3430 = ~n3427 & ~n3429;
  assign n3431 = ~A640  & A641 ;
  assign n3432 = A640  & ~A641 ;
  assign n3433 = A642  & ~n3432;
  assign n3434 = ~n3431 & n3433;
  assign n3435 = ~n3431 & ~n3432;
  assign n3436 = ~A642  & ~n3435;
  assign n3437 = ~n3434 & ~n3436;
  assign n3438 = ~n3430 & n3437;
  assign n3439 = n3430 & ~n3437;
  assign n3440 = ~n3438 & ~n3439;
  assign n3441 = A640  & A641 ;
  assign n3442 = A642  & ~n3435;
  assign n3443 = ~n3441 & ~n3442;
  assign n3444 = A637  & A638 ;
  assign n3445 = A639  & ~n3428;
  assign n3446 = ~n3444 & ~n3445;
  assign n3447 = ~n3443 & n3446;
  assign n3448 = n3443 & ~n3446;
  assign n3449 = ~n3447 & ~n3448;
  assign n3450 = ~n3430 & ~n3437;
  assign n3451 = ~n3449 & n3450;
  assign n3452 = ~n3443 & ~n3446;
  assign n3453 = ~n3451 & ~n3452;
  assign n3454 = ~n3447 & n3450;
  assign n3455 = ~n3448 & n3454;
  assign n3456 = ~n3449 & ~n3450;
  assign n3457 = ~n3455 & ~n3456;
  assign n3458 = ~n3453 & ~n3457;
  assign n3459 = ~n3440 & ~n3458;
  assign n3460 = ~A631  & A632 ;
  assign n3461 = A631  & ~A632 ;
  assign n3462 = A633  & ~n3461;
  assign n3463 = ~n3460 & n3462;
  assign n3464 = ~n3460 & ~n3461;
  assign n3465 = ~A633  & ~n3464;
  assign n3466 = ~n3463 & ~n3465;
  assign n3467 = ~A634  & A635 ;
  assign n3468 = A634  & ~A635 ;
  assign n3469 = A636  & ~n3468;
  assign n3470 = ~n3467 & n3469;
  assign n3471 = ~n3467 & ~n3468;
  assign n3472 = ~A636  & ~n3471;
  assign n3473 = ~n3470 & ~n3472;
  assign n3474 = ~n3466 & n3473;
  assign n3475 = n3466 & ~n3473;
  assign n3476 = ~n3474 & ~n3475;
  assign n3477 = A634  & A635 ;
  assign n3478 = A636  & ~n3471;
  assign n3479 = ~n3477 & ~n3478;
  assign n3480 = A631  & A632 ;
  assign n3481 = A633  & ~n3464;
  assign n3482 = ~n3480 & ~n3481;
  assign n3483 = ~n3479 & n3482;
  assign n3484 = n3479 & ~n3482;
  assign n3485 = ~n3483 & ~n3484;
  assign n3486 = ~n3466 & ~n3473;
  assign n3487 = ~n3485 & n3486;
  assign n3488 = ~n3479 & ~n3482;
  assign n3489 = ~n3487 & ~n3488;
  assign n3490 = ~n3483 & n3486;
  assign n3491 = ~n3484 & n3490;
  assign n3492 = ~n3485 & ~n3486;
  assign n3493 = ~n3491 & ~n3492;
  assign n3494 = ~n3489 & ~n3493;
  assign n3495 = ~n3476 & ~n3494;
  assign n3496 = ~n3459 & n3495;
  assign n3497 = n3459 & ~n3495;
  assign n3498 = ~n3496 & ~n3497;
  assign n3499 = ~n3423 & n3498;
  assign n3500 = n3423 & ~n3498;
  assign n3501 = ~n3499 & ~n3500;
  assign n3502 = ~A625  & A626 ;
  assign n3503 = A625  & ~A626 ;
  assign n3504 = A627  & ~n3503;
  assign n3505 = ~n3502 & n3504;
  assign n3506 = ~n3502 & ~n3503;
  assign n3507 = ~A627  & ~n3506;
  assign n3508 = ~n3505 & ~n3507;
  assign n3509 = ~A628  & A629 ;
  assign n3510 = A628  & ~A629 ;
  assign n3511 = A630  & ~n3510;
  assign n3512 = ~n3509 & n3511;
  assign n3513 = ~n3509 & ~n3510;
  assign n3514 = ~A630  & ~n3513;
  assign n3515 = ~n3512 & ~n3514;
  assign n3516 = ~n3508 & n3515;
  assign n3517 = n3508 & ~n3515;
  assign n3518 = ~n3516 & ~n3517;
  assign n3519 = A628  & A629 ;
  assign n3520 = A630  & ~n3513;
  assign n3521 = ~n3519 & ~n3520;
  assign n3522 = A625  & A626 ;
  assign n3523 = A627  & ~n3506;
  assign n3524 = ~n3522 & ~n3523;
  assign n3525 = ~n3521 & n3524;
  assign n3526 = n3521 & ~n3524;
  assign n3527 = ~n3525 & ~n3526;
  assign n3528 = ~n3508 & ~n3515;
  assign n3529 = ~n3527 & n3528;
  assign n3530 = ~n3521 & ~n3524;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = ~n3525 & n3528;
  assign n3533 = ~n3526 & n3532;
  assign n3534 = ~n3527 & ~n3528;
  assign n3535 = ~n3533 & ~n3534;
  assign n3536 = ~n3531 & ~n3535;
  assign n3537 = ~n3518 & ~n3536;
  assign n3538 = ~A619  & A620 ;
  assign n3539 = A619  & ~A620 ;
  assign n3540 = A621  & ~n3539;
  assign n3541 = ~n3538 & n3540;
  assign n3542 = ~n3538 & ~n3539;
  assign n3543 = ~A621  & ~n3542;
  assign n3544 = ~n3541 & ~n3543;
  assign n3545 = ~A622  & A623 ;
  assign n3546 = A622  & ~A623 ;
  assign n3547 = A624  & ~n3546;
  assign n3548 = ~n3545 & n3547;
  assign n3549 = ~n3545 & ~n3546;
  assign n3550 = ~A624  & ~n3549;
  assign n3551 = ~n3548 & ~n3550;
  assign n3552 = ~n3544 & n3551;
  assign n3553 = n3544 & ~n3551;
  assign n3554 = ~n3552 & ~n3553;
  assign n3555 = A622  & A623 ;
  assign n3556 = A624  & ~n3549;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = A619  & A620 ;
  assign n3559 = A621  & ~n3542;
  assign n3560 = ~n3558 & ~n3559;
  assign n3561 = ~n3557 & n3560;
  assign n3562 = n3557 & ~n3560;
  assign n3563 = ~n3561 & ~n3562;
  assign n3564 = ~n3544 & ~n3551;
  assign n3565 = ~n3563 & n3564;
  assign n3566 = ~n3557 & ~n3560;
  assign n3567 = ~n3565 & ~n3566;
  assign n3568 = ~n3561 & n3564;
  assign n3569 = ~n3562 & n3568;
  assign n3570 = ~n3563 & ~n3564;
  assign n3571 = ~n3569 & ~n3570;
  assign n3572 = ~n3567 & ~n3571;
  assign n3573 = ~n3554 & ~n3572;
  assign n3574 = ~n3537 & n3573;
  assign n3575 = n3537 & ~n3573;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = ~A613  & A614 ;
  assign n3578 = A613  & ~A614 ;
  assign n3579 = A615  & ~n3578;
  assign n3580 = ~n3577 & n3579;
  assign n3581 = ~n3577 & ~n3578;
  assign n3582 = ~A615  & ~n3581;
  assign n3583 = ~n3580 & ~n3582;
  assign n3584 = ~A616  & A617 ;
  assign n3585 = A616  & ~A617 ;
  assign n3586 = A618  & ~n3585;
  assign n3587 = ~n3584 & n3586;
  assign n3588 = ~n3584 & ~n3585;
  assign n3589 = ~A618  & ~n3588;
  assign n3590 = ~n3587 & ~n3589;
  assign n3591 = ~n3583 & n3590;
  assign n3592 = n3583 & ~n3590;
  assign n3593 = ~n3591 & ~n3592;
  assign n3594 = A616  & A617 ;
  assign n3595 = A618  & ~n3588;
  assign n3596 = ~n3594 & ~n3595;
  assign n3597 = A613  & A614 ;
  assign n3598 = A615  & ~n3581;
  assign n3599 = ~n3597 & ~n3598;
  assign n3600 = ~n3596 & n3599;
  assign n3601 = n3596 & ~n3599;
  assign n3602 = ~n3600 & ~n3601;
  assign n3603 = ~n3583 & ~n3590;
  assign n3604 = ~n3602 & n3603;
  assign n3605 = ~n3596 & ~n3599;
  assign n3606 = ~n3604 & ~n3605;
  assign n3607 = ~n3600 & n3603;
  assign n3608 = ~n3601 & n3607;
  assign n3609 = ~n3602 & ~n3603;
  assign n3610 = ~n3608 & ~n3609;
  assign n3611 = ~n3606 & ~n3610;
  assign n3612 = ~n3593 & ~n3611;
  assign n3613 = ~A607  & A608 ;
  assign n3614 = A607  & ~A608 ;
  assign n3615 = A609  & ~n3614;
  assign n3616 = ~n3613 & n3615;
  assign n3617 = ~n3613 & ~n3614;
  assign n3618 = ~A609  & ~n3617;
  assign n3619 = ~n3616 & ~n3618;
  assign n3620 = ~A610  & A611 ;
  assign n3621 = A610  & ~A611 ;
  assign n3622 = A612  & ~n3621;
  assign n3623 = ~n3620 & n3622;
  assign n3624 = ~n3620 & ~n3621;
  assign n3625 = ~A612  & ~n3624;
  assign n3626 = ~n3623 & ~n3625;
  assign n3627 = ~n3619 & n3626;
  assign n3628 = n3619 & ~n3626;
  assign n3629 = ~n3627 & ~n3628;
  assign n3630 = A610  & A611 ;
  assign n3631 = A612  & ~n3624;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = A607  & A608 ;
  assign n3634 = A609  & ~n3617;
  assign n3635 = ~n3633 & ~n3634;
  assign n3636 = ~n3632 & n3635;
  assign n3637 = n3632 & ~n3635;
  assign n3638 = ~n3636 & ~n3637;
  assign n3639 = ~n3619 & ~n3626;
  assign n3640 = ~n3638 & n3639;
  assign n3641 = ~n3632 & ~n3635;
  assign n3642 = ~n3640 & ~n3641;
  assign n3643 = ~n3636 & n3639;
  assign n3644 = ~n3637 & n3643;
  assign n3645 = ~n3638 & ~n3639;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = ~n3642 & ~n3646;
  assign n3648 = ~n3629 & ~n3647;
  assign n3649 = ~n3612 & n3648;
  assign n3650 = n3612 & ~n3648;
  assign n3651 = ~n3649 & ~n3650;
  assign n3652 = ~n3576 & n3651;
  assign n3653 = n3576 & ~n3651;
  assign n3654 = ~n3652 & ~n3653;
  assign n3655 = ~n3501 & n3654;
  assign n3656 = n3501 & ~n3654;
  assign n3657 = ~n3655 & ~n3656;
  assign n3658 = ~A601  & A602 ;
  assign n3659 = A601  & ~A602 ;
  assign n3660 = A603  & ~n3659;
  assign n3661 = ~n3658 & n3660;
  assign n3662 = ~n3658 & ~n3659;
  assign n3663 = ~A603  & ~n3662;
  assign n3664 = ~n3661 & ~n3663;
  assign n3665 = ~A604  & A605 ;
  assign n3666 = A604  & ~A605 ;
  assign n3667 = A606  & ~n3666;
  assign n3668 = ~n3665 & n3667;
  assign n3669 = ~n3665 & ~n3666;
  assign n3670 = ~A606  & ~n3669;
  assign n3671 = ~n3668 & ~n3670;
  assign n3672 = ~n3664 & n3671;
  assign n3673 = n3664 & ~n3671;
  assign n3674 = ~n3672 & ~n3673;
  assign n3675 = A604  & A605 ;
  assign n3676 = A606  & ~n3669;
  assign n3677 = ~n3675 & ~n3676;
  assign n3678 = A601  & A602 ;
  assign n3679 = A603  & ~n3662;
  assign n3680 = ~n3678 & ~n3679;
  assign n3681 = ~n3677 & n3680;
  assign n3682 = n3677 & ~n3680;
  assign n3683 = ~n3681 & ~n3682;
  assign n3684 = ~n3664 & ~n3671;
  assign n3685 = ~n3683 & n3684;
  assign n3686 = ~n3677 & ~n3680;
  assign n3687 = ~n3685 & ~n3686;
  assign n3688 = ~n3681 & n3684;
  assign n3689 = ~n3682 & n3688;
  assign n3690 = ~n3683 & ~n3684;
  assign n3691 = ~n3689 & ~n3690;
  assign n3692 = ~n3687 & ~n3691;
  assign n3693 = ~n3674 & ~n3692;
  assign n3694 = ~A595  & A596 ;
  assign n3695 = A595  & ~A596 ;
  assign n3696 = A597  & ~n3695;
  assign n3697 = ~n3694 & n3696;
  assign n3698 = ~n3694 & ~n3695;
  assign n3699 = ~A597  & ~n3698;
  assign n3700 = ~n3697 & ~n3699;
  assign n3701 = ~A598  & A599 ;
  assign n3702 = A598  & ~A599 ;
  assign n3703 = A600  & ~n3702;
  assign n3704 = ~n3701 & n3703;
  assign n3705 = ~n3701 & ~n3702;
  assign n3706 = ~A600  & ~n3705;
  assign n3707 = ~n3704 & ~n3706;
  assign n3708 = ~n3700 & n3707;
  assign n3709 = n3700 & ~n3707;
  assign n3710 = ~n3708 & ~n3709;
  assign n3711 = A598  & A599 ;
  assign n3712 = A600  & ~n3705;
  assign n3713 = ~n3711 & ~n3712;
  assign n3714 = A595  & A596 ;
  assign n3715 = A597  & ~n3698;
  assign n3716 = ~n3714 & ~n3715;
  assign n3717 = ~n3713 & n3716;
  assign n3718 = n3713 & ~n3716;
  assign n3719 = ~n3717 & ~n3718;
  assign n3720 = ~n3700 & ~n3707;
  assign n3721 = ~n3719 & n3720;
  assign n3722 = ~n3713 & ~n3716;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = ~n3717 & n3720;
  assign n3725 = ~n3718 & n3724;
  assign n3726 = ~n3719 & ~n3720;
  assign n3727 = ~n3725 & ~n3726;
  assign n3728 = ~n3723 & ~n3727;
  assign n3729 = ~n3710 & ~n3728;
  assign n3730 = ~n3693 & n3729;
  assign n3731 = n3693 & ~n3729;
  assign n3732 = ~n3730 & ~n3731;
  assign n3733 = ~A589  & A590 ;
  assign n3734 = A589  & ~A590 ;
  assign n3735 = A591  & ~n3734;
  assign n3736 = ~n3733 & n3735;
  assign n3737 = ~n3733 & ~n3734;
  assign n3738 = ~A591  & ~n3737;
  assign n3739 = ~n3736 & ~n3738;
  assign n3740 = ~A592  & A593 ;
  assign n3741 = A592  & ~A593 ;
  assign n3742 = A594  & ~n3741;
  assign n3743 = ~n3740 & n3742;
  assign n3744 = ~n3740 & ~n3741;
  assign n3745 = ~A594  & ~n3744;
  assign n3746 = ~n3743 & ~n3745;
  assign n3747 = ~n3739 & n3746;
  assign n3748 = n3739 & ~n3746;
  assign n3749 = ~n3747 & ~n3748;
  assign n3750 = A592  & A593 ;
  assign n3751 = A594  & ~n3744;
  assign n3752 = ~n3750 & ~n3751;
  assign n3753 = A589  & A590 ;
  assign n3754 = A591  & ~n3737;
  assign n3755 = ~n3753 & ~n3754;
  assign n3756 = ~n3752 & n3755;
  assign n3757 = n3752 & ~n3755;
  assign n3758 = ~n3756 & ~n3757;
  assign n3759 = ~n3739 & ~n3746;
  assign n3760 = ~n3758 & n3759;
  assign n3761 = ~n3752 & ~n3755;
  assign n3762 = ~n3760 & ~n3761;
  assign n3763 = ~n3756 & n3759;
  assign n3764 = ~n3757 & n3763;
  assign n3765 = ~n3758 & ~n3759;
  assign n3766 = ~n3764 & ~n3765;
  assign n3767 = ~n3762 & ~n3766;
  assign n3768 = ~n3749 & ~n3767;
  assign n3769 = ~A583  & A584 ;
  assign n3770 = A583  & ~A584 ;
  assign n3771 = A585  & ~n3770;
  assign n3772 = ~n3769 & n3771;
  assign n3773 = ~n3769 & ~n3770;
  assign n3774 = ~A585  & ~n3773;
  assign n3775 = ~n3772 & ~n3774;
  assign n3776 = ~A586  & A587 ;
  assign n3777 = A586  & ~A587 ;
  assign n3778 = A588  & ~n3777;
  assign n3779 = ~n3776 & n3778;
  assign n3780 = ~n3776 & ~n3777;
  assign n3781 = ~A588  & ~n3780;
  assign n3782 = ~n3779 & ~n3781;
  assign n3783 = ~n3775 & n3782;
  assign n3784 = n3775 & ~n3782;
  assign n3785 = ~n3783 & ~n3784;
  assign n3786 = A586  & A587 ;
  assign n3787 = A588  & ~n3780;
  assign n3788 = ~n3786 & ~n3787;
  assign n3789 = A583  & A584 ;
  assign n3790 = A585  & ~n3773;
  assign n3791 = ~n3789 & ~n3790;
  assign n3792 = ~n3788 & n3791;
  assign n3793 = n3788 & ~n3791;
  assign n3794 = ~n3792 & ~n3793;
  assign n3795 = ~n3775 & ~n3782;
  assign n3796 = ~n3794 & n3795;
  assign n3797 = ~n3788 & ~n3791;
  assign n3798 = ~n3796 & ~n3797;
  assign n3799 = ~n3792 & n3795;
  assign n3800 = ~n3793 & n3799;
  assign n3801 = ~n3794 & ~n3795;
  assign n3802 = ~n3800 & ~n3801;
  assign n3803 = ~n3798 & ~n3802;
  assign n3804 = ~n3785 & ~n3803;
  assign n3805 = ~n3768 & n3804;
  assign n3806 = n3768 & ~n3804;
  assign n3807 = ~n3805 & ~n3806;
  assign n3808 = ~n3732 & n3807;
  assign n3809 = n3732 & ~n3807;
  assign n3810 = ~n3808 & ~n3809;
  assign n3811 = ~A577  & A578 ;
  assign n3812 = A577  & ~A578 ;
  assign n3813 = A579  & ~n3812;
  assign n3814 = ~n3811 & n3813;
  assign n3815 = ~n3811 & ~n3812;
  assign n3816 = ~A579  & ~n3815;
  assign n3817 = ~n3814 & ~n3816;
  assign n3818 = ~A580  & A581 ;
  assign n3819 = A580  & ~A581 ;
  assign n3820 = A582  & ~n3819;
  assign n3821 = ~n3818 & n3820;
  assign n3822 = ~n3818 & ~n3819;
  assign n3823 = ~A582  & ~n3822;
  assign n3824 = ~n3821 & ~n3823;
  assign n3825 = ~n3817 & n3824;
  assign n3826 = n3817 & ~n3824;
  assign n3827 = ~n3825 & ~n3826;
  assign n3828 = A580  & A581 ;
  assign n3829 = A582  & ~n3822;
  assign n3830 = ~n3828 & ~n3829;
  assign n3831 = A577  & A578 ;
  assign n3832 = A579  & ~n3815;
  assign n3833 = ~n3831 & ~n3832;
  assign n3834 = ~n3830 & n3833;
  assign n3835 = n3830 & ~n3833;
  assign n3836 = ~n3834 & ~n3835;
  assign n3837 = ~n3817 & ~n3824;
  assign n3838 = ~n3836 & n3837;
  assign n3839 = ~n3830 & ~n3833;
  assign n3840 = ~n3838 & ~n3839;
  assign n3841 = ~n3834 & n3837;
  assign n3842 = ~n3835 & n3841;
  assign n3843 = ~n3836 & ~n3837;
  assign n3844 = ~n3842 & ~n3843;
  assign n3845 = ~n3840 & ~n3844;
  assign n3846 = ~n3827 & ~n3845;
  assign n3847 = ~A571  & A572 ;
  assign n3848 = A571  & ~A572 ;
  assign n3849 = A573  & ~n3848;
  assign n3850 = ~n3847 & n3849;
  assign n3851 = ~n3847 & ~n3848;
  assign n3852 = ~A573  & ~n3851;
  assign n3853 = ~n3850 & ~n3852;
  assign n3854 = ~A574  & A575 ;
  assign n3855 = A574  & ~A575 ;
  assign n3856 = A576  & ~n3855;
  assign n3857 = ~n3854 & n3856;
  assign n3858 = ~n3854 & ~n3855;
  assign n3859 = ~A576  & ~n3858;
  assign n3860 = ~n3857 & ~n3859;
  assign n3861 = ~n3853 & n3860;
  assign n3862 = n3853 & ~n3860;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = A574  & A575 ;
  assign n3865 = A576  & ~n3858;
  assign n3866 = ~n3864 & ~n3865;
  assign n3867 = A571  & A572 ;
  assign n3868 = A573  & ~n3851;
  assign n3869 = ~n3867 & ~n3868;
  assign n3870 = ~n3866 & n3869;
  assign n3871 = n3866 & ~n3869;
  assign n3872 = ~n3870 & ~n3871;
  assign n3873 = ~n3853 & ~n3860;
  assign n3874 = ~n3872 & n3873;
  assign n3875 = ~n3866 & ~n3869;
  assign n3876 = ~n3874 & ~n3875;
  assign n3877 = ~n3870 & n3873;
  assign n3878 = ~n3871 & n3877;
  assign n3879 = ~n3872 & ~n3873;
  assign n3880 = ~n3878 & ~n3879;
  assign n3881 = ~n3876 & ~n3880;
  assign n3882 = ~n3863 & ~n3881;
  assign n3883 = ~n3846 & n3882;
  assign n3884 = n3846 & ~n3882;
  assign n3885 = ~n3883 & ~n3884;
  assign n3886 = ~A565  & A566 ;
  assign n3887 = A565  & ~A566 ;
  assign n3888 = A567  & ~n3887;
  assign n3889 = ~n3886 & n3888;
  assign n3890 = ~n3886 & ~n3887;
  assign n3891 = ~A567  & ~n3890;
  assign n3892 = ~n3889 & ~n3891;
  assign n3893 = ~A568  & A569 ;
  assign n3894 = A568  & ~A569 ;
  assign n3895 = A570  & ~n3894;
  assign n3896 = ~n3893 & n3895;
  assign n3897 = ~n3893 & ~n3894;
  assign n3898 = ~A570  & ~n3897;
  assign n3899 = ~n3896 & ~n3898;
  assign n3900 = ~n3892 & n3899;
  assign n3901 = n3892 & ~n3899;
  assign n3902 = ~n3900 & ~n3901;
  assign n3903 = A568  & A569 ;
  assign n3904 = A570  & ~n3897;
  assign n3905 = ~n3903 & ~n3904;
  assign n3906 = A565  & A566 ;
  assign n3907 = A567  & ~n3890;
  assign n3908 = ~n3906 & ~n3907;
  assign n3909 = ~n3905 & n3908;
  assign n3910 = n3905 & ~n3908;
  assign n3911 = ~n3909 & ~n3910;
  assign n3912 = ~n3892 & ~n3899;
  assign n3913 = ~n3911 & n3912;
  assign n3914 = ~n3905 & ~n3908;
  assign n3915 = ~n3913 & ~n3914;
  assign n3916 = ~n3909 & n3912;
  assign n3917 = ~n3910 & n3916;
  assign n3918 = ~n3911 & ~n3912;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = ~n3915 & ~n3919;
  assign n3921 = ~n3902 & ~n3920;
  assign n3922 = ~A559  & A560 ;
  assign n3923 = A559  & ~A560 ;
  assign n3924 = A561  & ~n3923;
  assign n3925 = ~n3922 & n3924;
  assign n3926 = ~n3922 & ~n3923;
  assign n3927 = ~A561  & ~n3926;
  assign n3928 = ~n3925 & ~n3927;
  assign n3929 = ~A562  & A563 ;
  assign n3930 = A562  & ~A563 ;
  assign n3931 = A564  & ~n3930;
  assign n3932 = ~n3929 & n3931;
  assign n3933 = ~n3929 & ~n3930;
  assign n3934 = ~A564  & ~n3933;
  assign n3935 = ~n3932 & ~n3934;
  assign n3936 = ~n3928 & n3935;
  assign n3937 = n3928 & ~n3935;
  assign n3938 = ~n3936 & ~n3937;
  assign n3939 = A562  & A563 ;
  assign n3940 = A564  & ~n3933;
  assign n3941 = ~n3939 & ~n3940;
  assign n3942 = A559  & A560 ;
  assign n3943 = A561  & ~n3926;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = ~n3941 & n3944;
  assign n3946 = n3941 & ~n3944;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = ~n3928 & ~n3935;
  assign n3949 = ~n3947 & n3948;
  assign n3950 = ~n3941 & ~n3944;
  assign n3951 = ~n3949 & ~n3950;
  assign n3952 = ~n3945 & n3948;
  assign n3953 = ~n3946 & n3952;
  assign n3954 = ~n3947 & ~n3948;
  assign n3955 = ~n3953 & ~n3954;
  assign n3956 = ~n3951 & ~n3955;
  assign n3957 = ~n3938 & ~n3956;
  assign n3958 = ~n3921 & n3957;
  assign n3959 = n3921 & ~n3957;
  assign n3960 = ~n3958 & ~n3959;
  assign n3961 = ~n3885 & n3960;
  assign n3962 = n3885 & ~n3960;
  assign n3963 = ~n3961 & ~n3962;
  assign n3964 = ~n3810 & n3963;
  assign n3965 = n3810 & ~n3963;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = ~n3657 & n3966;
  assign n3968 = n3657 & ~n3966;
  assign n3969 = ~n3967 & ~n3968;
  assign n3970 = ~n3348 & n3969;
  assign n3971 = n3348 & ~n3969;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = ~n2712 & n2715;
  assign n3974 = n2712 & ~n2715;
  assign n3975 = ~n3973 & ~n3974;
  assign n3976 = ~n3972 & ~n3975;
  assign n3977 = ~n2727 & n3976;
  assign n3978 = ~n2722 & n3977;
  assign n3979 = ~n2722 & ~n2727;
  assign n3980 = ~n3976 & ~n3979;
  assign n3981 = ~n3978 & ~n3980;
  assign n3982 = ~n3785 & ~n3798;
  assign n3983 = ~n3802 & ~n3982;
  assign n3984 = ~n3749 & ~n3785;
  assign n3985 = ~n3767 & n3984;
  assign n3986 = ~n3803 & n3985;
  assign n3987 = ~n3749 & ~n3762;
  assign n3988 = ~n3766 & ~n3987;
  assign n3989 = ~n3986 & n3988;
  assign n3990 = n3986 & ~n3988;
  assign n3991 = ~n3989 & ~n3990;
  assign n3992 = ~n3983 & ~n3991;
  assign n3993 = ~n3986 & ~n3988;
  assign n3994 = ~n3766 & n3984;
  assign n3995 = ~n3767 & n3994;
  assign n3996 = ~n3803 & ~n3987;
  assign n3997 = n3995 & n3996;
  assign n3998 = ~n3993 & ~n3997;
  assign n3999 = n3983 & ~n3998;
  assign n4000 = ~n3992 & ~n3999;
  assign n4001 = ~n3710 & ~n3723;
  assign n4002 = ~n3727 & ~n4001;
  assign n4003 = ~n3674 & ~n3710;
  assign n4004 = ~n3692 & n4003;
  assign n4005 = ~n3728 & n4004;
  assign n4006 = ~n3674 & ~n3687;
  assign n4007 = ~n3691 & ~n4006;
  assign n4008 = ~n4005 & ~n4007;
  assign n4009 = ~n3691 & n4003;
  assign n4010 = ~n3692 & n4009;
  assign n4011 = ~n3728 & ~n4006;
  assign n4012 = n4010 & n4011;
  assign n4013 = ~n4008 & ~n4012;
  assign n4014 = n4002 & ~n4013;
  assign n4015 = ~n4005 & n4007;
  assign n4016 = n4005 & ~n4007;
  assign n4017 = ~n4015 & ~n4016;
  assign n4018 = ~n4002 & ~n4017;
  assign n4019 = ~n3732 & ~n3807;
  assign n4020 = ~n4018 & ~n4019;
  assign n4021 = ~n4014 & n4020;
  assign n4022 = ~n4014 & ~n4018;
  assign n4023 = n4019 & ~n4022;
  assign n4024 = ~n4021 & ~n4023;
  assign n4025 = ~n4000 & ~n4024;
  assign n4026 = ~n4018 & n4019;
  assign n4027 = ~n4014 & n4026;
  assign n4028 = ~n4019 & ~n4022;
  assign n4029 = ~n4027 & ~n4028;
  assign n4030 = n4000 & ~n4029;
  assign n4031 = ~n3810 & ~n3963;
  assign n4032 = ~n4030 & n4031;
  assign n4033 = ~n4025 & n4032;
  assign n4034 = ~n4025 & ~n4030;
  assign n4035 = ~n4031 & ~n4034;
  assign n4036 = ~n4033 & ~n4035;
  assign n4037 = ~n3863 & ~n3876;
  assign n4038 = ~n3880 & ~n4037;
  assign n4039 = ~n3827 & ~n3863;
  assign n4040 = ~n3845 & n4039;
  assign n4041 = ~n3881 & n4040;
  assign n4042 = ~n3827 & ~n3840;
  assign n4043 = ~n3844 & ~n4042;
  assign n4044 = ~n4041 & ~n4043;
  assign n4045 = ~n3844 & n4039;
  assign n4046 = ~n3845 & n4045;
  assign n4047 = ~n3881 & ~n4042;
  assign n4048 = n4046 & n4047;
  assign n4049 = ~n4044 & ~n4048;
  assign n4050 = n4038 & ~n4049;
  assign n4051 = ~n4041 & n4043;
  assign n4052 = n4041 & ~n4043;
  assign n4053 = ~n4051 & ~n4052;
  assign n4054 = ~n4038 & ~n4053;
  assign n4055 = ~n3885 & ~n3960;
  assign n4056 = ~n4054 & n4055;
  assign n4057 = ~n4050 & n4056;
  assign n4058 = ~n4050 & ~n4054;
  assign n4059 = ~n4055 & ~n4058;
  assign n4060 = ~n4057 & ~n4059;
  assign n4061 = ~n3938 & ~n3951;
  assign n4062 = ~n3955 & ~n4061;
  assign n4063 = ~n3902 & ~n3938;
  assign n4064 = ~n3920 & n4063;
  assign n4065 = ~n3956 & n4064;
  assign n4066 = ~n3902 & ~n3915;
  assign n4067 = ~n3919 & ~n4066;
  assign n4068 = ~n4065 & n4067;
  assign n4069 = n4065 & ~n4067;
  assign n4070 = ~n4068 & ~n4069;
  assign n4071 = ~n4062 & ~n4070;
  assign n4072 = ~n4065 & ~n4067;
  assign n4073 = ~n3919 & n4063;
  assign n4074 = ~n3920 & n4073;
  assign n4075 = ~n3956 & ~n4066;
  assign n4076 = n4074 & n4075;
  assign n4077 = ~n4072 & ~n4076;
  assign n4078 = n4062 & ~n4077;
  assign n4079 = ~n4071 & ~n4078;
  assign n4080 = ~n4060 & n4079;
  assign n4081 = ~n4054 & ~n4055;
  assign n4082 = ~n4050 & n4081;
  assign n4083 = n4055 & ~n4058;
  assign n4084 = ~n4082 & ~n4083;
  assign n4085 = ~n4079 & ~n4084;
  assign n4086 = ~n4080 & ~n4085;
  assign n4087 = ~n4036 & n4086;
  assign n4088 = ~n4030 & ~n4031;
  assign n4089 = ~n4025 & n4088;
  assign n4090 = n4031 & ~n4034;
  assign n4091 = ~n4089 & ~n4090;
  assign n4092 = ~n4086 & ~n4091;
  assign n4093 = ~n4087 & ~n4092;
  assign n4094 = ~n3554 & ~n3567;
  assign n4095 = ~n3571 & ~n4094;
  assign n4096 = ~n3518 & ~n3554;
  assign n4097 = ~n3536 & n4096;
  assign n4098 = ~n3572 & n4097;
  assign n4099 = ~n3518 & ~n3531;
  assign n4100 = ~n3535 & ~n4099;
  assign n4101 = ~n4098 & ~n4100;
  assign n4102 = ~n3535 & n4096;
  assign n4103 = ~n3536 & n4102;
  assign n4104 = ~n3572 & ~n4099;
  assign n4105 = n4103 & n4104;
  assign n4106 = ~n4101 & ~n4105;
  assign n4107 = n4095 & ~n4106;
  assign n4108 = ~n4098 & n4100;
  assign n4109 = n4098 & ~n4100;
  assign n4110 = ~n4108 & ~n4109;
  assign n4111 = ~n4095 & ~n4110;
  assign n4112 = ~n3576 & ~n3651;
  assign n4113 = ~n4111 & n4112;
  assign n4114 = ~n4107 & n4113;
  assign n4115 = ~n4107 & ~n4111;
  assign n4116 = ~n4112 & ~n4115;
  assign n4117 = ~n4114 & ~n4116;
  assign n4118 = ~n3629 & ~n3642;
  assign n4119 = ~n3646 & ~n4118;
  assign n4120 = ~n3593 & ~n3629;
  assign n4121 = ~n3611 & n4120;
  assign n4122 = ~n3647 & n4121;
  assign n4123 = ~n3593 & ~n3606;
  assign n4124 = ~n3610 & ~n4123;
  assign n4125 = ~n4122 & n4124;
  assign n4126 = n4122 & ~n4124;
  assign n4127 = ~n4125 & ~n4126;
  assign n4128 = ~n4119 & ~n4127;
  assign n4129 = ~n4122 & ~n4124;
  assign n4130 = ~n3610 & n4120;
  assign n4131 = ~n3611 & n4130;
  assign n4132 = ~n3647 & ~n4123;
  assign n4133 = n4131 & n4132;
  assign n4134 = ~n4129 & ~n4133;
  assign n4135 = n4119 & ~n4134;
  assign n4136 = ~n4128 & ~n4135;
  assign n4137 = ~n4117 & n4136;
  assign n4138 = ~n4111 & ~n4112;
  assign n4139 = ~n4107 & n4138;
  assign n4140 = n4112 & ~n4115;
  assign n4141 = ~n4139 & ~n4140;
  assign n4142 = ~n4136 & ~n4141;
  assign n4143 = ~n4137 & ~n4142;
  assign n4144 = ~n3476 & ~n3489;
  assign n4145 = ~n3493 & ~n4144;
  assign n4146 = ~n3440 & ~n3476;
  assign n4147 = ~n3458 & n4146;
  assign n4148 = ~n3494 & n4147;
  assign n4149 = ~n3440 & ~n3453;
  assign n4150 = ~n3457 & ~n4149;
  assign n4151 = ~n4148 & n4150;
  assign n4152 = n4148 & ~n4150;
  assign n4153 = ~n4151 & ~n4152;
  assign n4154 = ~n4145 & ~n4153;
  assign n4155 = ~n4148 & ~n4150;
  assign n4156 = ~n3457 & n4146;
  assign n4157 = ~n3458 & n4156;
  assign n4158 = ~n3494 & ~n4149;
  assign n4159 = n4157 & n4158;
  assign n4160 = ~n4155 & ~n4159;
  assign n4161 = n4145 & ~n4160;
  assign n4162 = ~n4154 & ~n4161;
  assign n4163 = ~n3401 & ~n3414;
  assign n4164 = ~n3418 & ~n4163;
  assign n4165 = ~n3365 & ~n3401;
  assign n4166 = ~n3383 & n4165;
  assign n4167 = ~n3419 & n4166;
  assign n4168 = ~n3365 & ~n3378;
  assign n4169 = ~n3382 & ~n4168;
  assign n4170 = ~n4167 & ~n4169;
  assign n4171 = ~n3382 & n4165;
  assign n4172 = ~n3383 & n4171;
  assign n4173 = ~n3419 & ~n4168;
  assign n4174 = n4172 & n4173;
  assign n4175 = ~n4170 & ~n4174;
  assign n4176 = n4164 & ~n4175;
  assign n4177 = ~n4167 & n4169;
  assign n4178 = n4167 & ~n4169;
  assign n4179 = ~n4177 & ~n4178;
  assign n4180 = ~n4164 & ~n4179;
  assign n4181 = ~n3423 & ~n3498;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = ~n4176 & n4182;
  assign n4184 = ~n4176 & ~n4180;
  assign n4185 = n4181 & ~n4184;
  assign n4186 = ~n4183 & ~n4185;
  assign n4187 = ~n4162 & ~n4186;
  assign n4188 = ~n4180 & n4181;
  assign n4189 = ~n4176 & n4188;
  assign n4190 = ~n4181 & ~n4184;
  assign n4191 = ~n4189 & ~n4190;
  assign n4192 = n4162 & ~n4191;
  assign n4193 = ~n3501 & ~n3654;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = ~n4187 & n4194;
  assign n4196 = ~n4187 & ~n4192;
  assign n4197 = n4193 & ~n4196;
  assign n4198 = ~n4195 & ~n4197;
  assign n4199 = ~n4143 & ~n4198;
  assign n4200 = ~n4192 & n4193;
  assign n4201 = ~n4187 & n4200;
  assign n4202 = ~n4193 & ~n4196;
  assign n4203 = ~n4201 & ~n4202;
  assign n4204 = n4143 & ~n4203;
  assign n4205 = ~n3657 & ~n3966;
  assign n4206 = ~n4204 & ~n4205;
  assign n4207 = ~n4199 & n4206;
  assign n4208 = ~n4199 & ~n4204;
  assign n4209 = n4205 & ~n4208;
  assign n4210 = ~n4207 & ~n4209;
  assign n4211 = ~n4093 & ~n4210;
  assign n4212 = ~n4204 & n4205;
  assign n4213 = ~n4199 & n4212;
  assign n4214 = ~n4205 & ~n4208;
  assign n4215 = ~n4213 & ~n4214;
  assign n4216 = n4093 & ~n4215;
  assign n4217 = ~n3348 & ~n3969;
  assign n4218 = ~n4216 & n4217;
  assign n4219 = ~n4211 & n4218;
  assign n4220 = ~n4211 & ~n4216;
  assign n4221 = ~n4217 & ~n4220;
  assign n4222 = ~n4219 & ~n4221;
  assign n4223 = ~n3242 & ~n3255;
  assign n4224 = ~n3259 & ~n4223;
  assign n4225 = ~n3206 & ~n3242;
  assign n4226 = ~n3224 & n4225;
  assign n4227 = ~n3260 & n4226;
  assign n4228 = ~n3206 & ~n3219;
  assign n4229 = ~n3223 & ~n4228;
  assign n4230 = ~n4227 & ~n4229;
  assign n4231 = ~n3223 & n4225;
  assign n4232 = ~n3224 & n4231;
  assign n4233 = ~n3260 & ~n4228;
  assign n4234 = n4232 & n4233;
  assign n4235 = ~n4230 & ~n4234;
  assign n4236 = n4224 & ~n4235;
  assign n4237 = ~n4227 & n4229;
  assign n4238 = n4227 & ~n4229;
  assign n4239 = ~n4237 & ~n4238;
  assign n4240 = ~n4224 & ~n4239;
  assign n4241 = ~n3264 & ~n3339;
  assign n4242 = ~n4240 & n4241;
  assign n4243 = ~n4236 & n4242;
  assign n4244 = ~n4236 & ~n4240;
  assign n4245 = ~n4241 & ~n4244;
  assign n4246 = ~n4243 & ~n4245;
  assign n4247 = ~n3317 & ~n3330;
  assign n4248 = ~n3334 & ~n4247;
  assign n4249 = ~n3281 & ~n3317;
  assign n4250 = ~n3299 & n4249;
  assign n4251 = ~n3335 & n4250;
  assign n4252 = ~n3281 & ~n3294;
  assign n4253 = ~n3298 & ~n4252;
  assign n4254 = ~n4251 & n4253;
  assign n4255 = n4251 & ~n4253;
  assign n4256 = ~n4254 & ~n4255;
  assign n4257 = ~n4248 & ~n4256;
  assign n4258 = ~n4251 & ~n4253;
  assign n4259 = ~n3298 & n4249;
  assign n4260 = ~n3299 & n4259;
  assign n4261 = ~n3335 & ~n4252;
  assign n4262 = n4260 & n4261;
  assign n4263 = ~n4258 & ~n4262;
  assign n4264 = n4248 & ~n4263;
  assign n4265 = ~n4257 & ~n4264;
  assign n4266 = ~n4246 & n4265;
  assign n4267 = ~n4240 & ~n4241;
  assign n4268 = ~n4236 & n4267;
  assign n4269 = n4241 & ~n4244;
  assign n4270 = ~n4268 & ~n4269;
  assign n4271 = ~n4265 & ~n4270;
  assign n4272 = ~n4266 & ~n4271;
  assign n4273 = ~n3164 & ~n3177;
  assign n4274 = ~n3181 & ~n4273;
  assign n4275 = ~n3128 & ~n3164;
  assign n4276 = ~n3146 & n4275;
  assign n4277 = ~n3182 & n4276;
  assign n4278 = ~n3128 & ~n3141;
  assign n4279 = ~n3145 & ~n4278;
  assign n4280 = ~n4277 & n4279;
  assign n4281 = n4277 & ~n4279;
  assign n4282 = ~n4280 & ~n4281;
  assign n4283 = ~n4274 & ~n4282;
  assign n4284 = ~n4277 & ~n4279;
  assign n4285 = ~n3145 & n4275;
  assign n4286 = ~n3146 & n4285;
  assign n4287 = ~n3182 & ~n4278;
  assign n4288 = n4286 & n4287;
  assign n4289 = ~n4284 & ~n4288;
  assign n4290 = n4274 & ~n4289;
  assign n4291 = ~n4283 & ~n4290;
  assign n4292 = ~n3089 & ~n3102;
  assign n4293 = ~n3106 & ~n4292;
  assign n4294 = ~n3053 & ~n3089;
  assign n4295 = ~n3071 & n4294;
  assign n4296 = ~n3107 & n4295;
  assign n4297 = ~n3053 & ~n3066;
  assign n4298 = ~n3070 & ~n4297;
  assign n4299 = ~n4296 & ~n4298;
  assign n4300 = ~n3070 & n4294;
  assign n4301 = ~n3071 & n4300;
  assign n4302 = ~n3107 & ~n4297;
  assign n4303 = n4301 & n4302;
  assign n4304 = ~n4299 & ~n4303;
  assign n4305 = n4293 & ~n4304;
  assign n4306 = ~n4296 & n4298;
  assign n4307 = n4296 & ~n4298;
  assign n4308 = ~n4306 & ~n4307;
  assign n4309 = ~n4293 & ~n4308;
  assign n4310 = ~n3111 & ~n3186;
  assign n4311 = ~n4309 & ~n4310;
  assign n4312 = ~n4305 & n4311;
  assign n4313 = ~n4305 & ~n4309;
  assign n4314 = n4310 & ~n4313;
  assign n4315 = ~n4312 & ~n4314;
  assign n4316 = ~n4291 & ~n4315;
  assign n4317 = ~n4309 & n4310;
  assign n4318 = ~n4305 & n4317;
  assign n4319 = ~n4310 & ~n4313;
  assign n4320 = ~n4318 & ~n4319;
  assign n4321 = n4291 & ~n4320;
  assign n4322 = ~n3189 & ~n3342;
  assign n4323 = ~n4321 & ~n4322;
  assign n4324 = ~n4316 & n4323;
  assign n4325 = ~n4316 & ~n4321;
  assign n4326 = n4322 & ~n4325;
  assign n4327 = ~n4324 & ~n4326;
  assign n4328 = ~n4272 & ~n4327;
  assign n4329 = ~n4321 & n4322;
  assign n4330 = ~n4316 & n4329;
  assign n4331 = ~n4322 & ~n4325;
  assign n4332 = ~n4330 & ~n4331;
  assign n4333 = n4272 & ~n4332;
  assign n4334 = ~n3036 & ~n3345;
  assign n4335 = ~n4333 & n4334;
  assign n4336 = ~n4328 & n4335;
  assign n4337 = ~n4328 & ~n4333;
  assign n4338 = ~n4334 & ~n4337;
  assign n4339 = ~n4336 & ~n4338;
  assign n4340 = ~n3008 & ~n3021;
  assign n4341 = ~n3025 & ~n4340;
  assign n4342 = ~n2972 & ~n3008;
  assign n4343 = ~n2990 & n4342;
  assign n4344 = ~n3026 & n4343;
  assign n4345 = ~n2972 & ~n2985;
  assign n4346 = ~n2989 & ~n4345;
  assign n4347 = ~n4344 & n4346;
  assign n4348 = n4344 & ~n4346;
  assign n4349 = ~n4347 & ~n4348;
  assign n4350 = ~n4341 & ~n4349;
  assign n4351 = ~n4344 & ~n4346;
  assign n4352 = ~n2989 & n4342;
  assign n4353 = ~n2990 & n4352;
  assign n4354 = ~n3026 & ~n4345;
  assign n4355 = n4353 & n4354;
  assign n4356 = ~n4351 & ~n4355;
  assign n4357 = n4341 & ~n4356;
  assign n4358 = ~n4350 & ~n4357;
  assign n4359 = ~n2933 & ~n2946;
  assign n4360 = ~n2950 & ~n4359;
  assign n4361 = ~n2897 & ~n2933;
  assign n4362 = ~n2915 & n4361;
  assign n4363 = ~n2951 & n4362;
  assign n4364 = ~n2897 & ~n2910;
  assign n4365 = ~n2914 & ~n4364;
  assign n4366 = ~n4363 & ~n4365;
  assign n4367 = ~n2914 & n4361;
  assign n4368 = ~n2915 & n4367;
  assign n4369 = ~n2951 & ~n4364;
  assign n4370 = n4368 & n4369;
  assign n4371 = ~n4366 & ~n4370;
  assign n4372 = n4360 & ~n4371;
  assign n4373 = ~n4363 & n4365;
  assign n4374 = n4363 & ~n4365;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = ~n4360 & ~n4375;
  assign n4377 = ~n2955 & ~n3030;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = ~n4372 & n4378;
  assign n4380 = ~n4372 & ~n4376;
  assign n4381 = n4377 & ~n4380;
  assign n4382 = ~n4379 & ~n4381;
  assign n4383 = ~n4358 & ~n4382;
  assign n4384 = ~n4376 & n4377;
  assign n4385 = ~n4372 & n4384;
  assign n4386 = ~n4377 & ~n4380;
  assign n4387 = ~n4385 & ~n4386;
  assign n4388 = n4358 & ~n4387;
  assign n4389 = ~n2880 & ~n3033;
  assign n4390 = ~n4388 & n4389;
  assign n4391 = ~n4383 & n4390;
  assign n4392 = ~n4383 & ~n4388;
  assign n4393 = ~n4389 & ~n4392;
  assign n4394 = ~n4391 & ~n4393;
  assign n4395 = ~n2855 & ~n2868;
  assign n4396 = ~n2872 & ~n4395;
  assign n4397 = ~n2819 & ~n2855;
  assign n4398 = ~n2837 & n4397;
  assign n4399 = ~n2873 & n4398;
  assign n4400 = ~n2819 & ~n2832;
  assign n4401 = ~n2836 & ~n4400;
  assign n4402 = ~n4399 & ~n4401;
  assign n4403 = ~n2836 & n4397;
  assign n4404 = ~n2837 & n4403;
  assign n4405 = ~n2873 & ~n4400;
  assign n4406 = n4404 & n4405;
  assign n4407 = ~n4402 & ~n4406;
  assign n4408 = n4396 & ~n4407;
  assign n4409 = ~n4399 & n4401;
  assign n4410 = n4399 & ~n4401;
  assign n4411 = ~n4409 & ~n4410;
  assign n4412 = ~n4396 & ~n4411;
  assign n4413 = ~n2802 & ~n2877;
  assign n4414 = ~n4412 & n4413;
  assign n4415 = ~n4408 & n4414;
  assign n4416 = ~n4408 & ~n4412;
  assign n4417 = ~n4413 & ~n4416;
  assign n4418 = ~n4415 & ~n4417;
  assign n4419 = ~n2780 & ~n2797;
  assign n4420 = ~n2794 & ~n4419;
  assign n4421 = ~n2744 & ~n2780;
  assign n4422 = ~n2762 & n4421;
  assign n4423 = ~n2798 & n4422;
  assign n4424 = ~n2744 & ~n2757;
  assign n4425 = ~n2761 & ~n4424;
  assign n4426 = ~n4423 & n4425;
  assign n4427 = n4423 & ~n4425;
  assign n4428 = ~n4426 & ~n4427;
  assign n4429 = ~n4420 & ~n4428;
  assign n4430 = ~n4423 & ~n4425;
  assign n4431 = ~n2761 & n4421;
  assign n4432 = ~n2762 & n4431;
  assign n4433 = ~n2798 & ~n4424;
  assign n4434 = n4432 & n4433;
  assign n4435 = ~n4430 & ~n4434;
  assign n4436 = n4420 & ~n4435;
  assign n4437 = ~n4429 & ~n4436;
  assign n4438 = ~n4418 & n4437;
  assign n4439 = ~n4412 & ~n4413;
  assign n4440 = ~n4408 & n4439;
  assign n4441 = n4413 & ~n4416;
  assign n4442 = ~n4440 & ~n4441;
  assign n4443 = ~n4437 & ~n4442;
  assign n4444 = ~n4438 & ~n4443;
  assign n4445 = ~n4394 & n4444;
  assign n4446 = ~n4388 & ~n4389;
  assign n4447 = ~n4383 & n4446;
  assign n4448 = n4389 & ~n4392;
  assign n4449 = ~n4447 & ~n4448;
  assign n4450 = ~n4444 & ~n4449;
  assign n4451 = ~n4445 & ~n4450;
  assign n4452 = ~n4339 & n4451;
  assign n4453 = ~n4333 & ~n4334;
  assign n4454 = ~n4328 & n4453;
  assign n4455 = n4334 & ~n4337;
  assign n4456 = ~n4454 & ~n4455;
  assign n4457 = ~n4451 & ~n4456;
  assign n4458 = ~n4452 & ~n4457;
  assign n4459 = ~n4222 & n4458;
  assign n4460 = ~n4216 & ~n4217;
  assign n4461 = ~n4211 & n4460;
  assign n4462 = n4217 & ~n4220;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = ~n4458 & ~n4463;
  assign n4465 = ~n4459 & ~n4464;
  assign n4466 = ~n3981 & n4465;
  assign n4467 = ~n2727 & ~n3976;
  assign n4468 = ~n2722 & n4467;
  assign n4469 = n3976 & ~n3979;
  assign n4470 = ~n4468 & ~n4469;
  assign n4471 = ~n4465 & ~n4470;
  assign n4472 = ~n4466 & ~n4471;
  assign n4473 = A970  & A971 ;
  assign n4474 = A970  & ~A971 ;
  assign n4475 = ~A970  & A971 ;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = A972  & ~n4476;
  assign n4478 = ~n4473 & ~n4477;
  assign n4479 = A967  & A968 ;
  assign n4480 = A967  & ~A968 ;
  assign n4481 = ~A967  & A968 ;
  assign n4482 = ~n4480 & ~n4481;
  assign n4483 = A969  & ~n4482;
  assign n4484 = ~n4479 & ~n4483;
  assign n4485 = n4478 & ~n4484;
  assign n4486 = ~n4478 & n4484;
  assign n4487 = A969  & ~n4480;
  assign n4488 = ~n4481 & n4487;
  assign n4489 = ~A969  & ~n4482;
  assign n4490 = ~n4488 & ~n4489;
  assign n4491 = A972  & ~n4474;
  assign n4492 = ~n4475 & n4491;
  assign n4493 = ~A972  & ~n4476;
  assign n4494 = ~n4492 & ~n4493;
  assign n4495 = ~n4490 & ~n4494;
  assign n4496 = ~n4486 & n4495;
  assign n4497 = ~n4485 & n4496;
  assign n4498 = ~n4485 & ~n4486;
  assign n4499 = ~n4495 & ~n4498;
  assign n4500 = ~n4497 & ~n4499;
  assign n4501 = ~n4490 & n4494;
  assign n4502 = n4490 & ~n4494;
  assign n4503 = ~n4501 & ~n4502;
  assign n4504 = n4495 & ~n4498;
  assign n4505 = ~n4478 & ~n4484;
  assign n4506 = ~n4504 & ~n4505;
  assign n4507 = ~n4503 & ~n4506;
  assign n4508 = ~n4500 & ~n4507;
  assign n4509 = ~n4500 & ~n4506;
  assign n4510 = A976  & A977 ;
  assign n4511 = A976  & ~A977 ;
  assign n4512 = ~A976  & A977 ;
  assign n4513 = ~n4511 & ~n4512;
  assign n4514 = A978  & ~n4513;
  assign n4515 = ~n4510 & ~n4514;
  assign n4516 = A973  & A974 ;
  assign n4517 = A973  & ~A974 ;
  assign n4518 = ~A973  & A974 ;
  assign n4519 = ~n4517 & ~n4518;
  assign n4520 = A975  & ~n4519;
  assign n4521 = ~n4516 & ~n4520;
  assign n4522 = ~n4515 & n4521;
  assign n4523 = n4515 & ~n4521;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = A975  & ~n4517;
  assign n4526 = ~n4518 & n4525;
  assign n4527 = ~A975  & ~n4519;
  assign n4528 = ~n4526 & ~n4527;
  assign n4529 = A978  & ~n4511;
  assign n4530 = ~n4512 & n4529;
  assign n4531 = ~A978  & ~n4513;
  assign n4532 = ~n4530 & ~n4531;
  assign n4533 = ~n4528 & ~n4532;
  assign n4534 = ~n4524 & n4533;
  assign n4535 = ~n4515 & ~n4521;
  assign n4536 = ~n4534 & ~n4535;
  assign n4537 = ~n4522 & n4533;
  assign n4538 = ~n4523 & n4537;
  assign n4539 = ~n4524 & ~n4533;
  assign n4540 = ~n4538 & ~n4539;
  assign n4541 = ~n4536 & ~n4540;
  assign n4542 = ~n4528 & n4532;
  assign n4543 = n4528 & ~n4532;
  assign n4544 = ~n4542 & ~n4543;
  assign n4545 = ~n4503 & ~n4544;
  assign n4546 = ~n4541 & n4545;
  assign n4547 = ~n4509 & n4546;
  assign n4548 = ~n4536 & ~n4544;
  assign n4549 = ~n4540 & ~n4548;
  assign n4550 = ~n4547 & n4549;
  assign n4551 = n4547 & ~n4549;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = ~n4508 & ~n4552;
  assign n4554 = ~n4547 & ~n4549;
  assign n4555 = ~n4540 & n4545;
  assign n4556 = ~n4541 & n4555;
  assign n4557 = ~n4509 & ~n4548;
  assign n4558 = n4556 & n4557;
  assign n4559 = ~n4554 & ~n4558;
  assign n4560 = n4508 & ~n4559;
  assign n4561 = ~n4553 & ~n4560;
  assign n4562 = A982  & A983 ;
  assign n4563 = A982  & ~A983 ;
  assign n4564 = ~A982  & A983 ;
  assign n4565 = ~n4563 & ~n4564;
  assign n4566 = A984  & ~n4565;
  assign n4567 = ~n4562 & ~n4566;
  assign n4568 = A979  & A980 ;
  assign n4569 = A979  & ~A980 ;
  assign n4570 = ~A979  & A980 ;
  assign n4571 = ~n4569 & ~n4570;
  assign n4572 = A981  & ~n4571;
  assign n4573 = ~n4568 & ~n4572;
  assign n4574 = n4567 & ~n4573;
  assign n4575 = ~n4567 & n4573;
  assign n4576 = A981  & ~n4569;
  assign n4577 = ~n4570 & n4576;
  assign n4578 = ~A981  & ~n4571;
  assign n4579 = ~n4577 & ~n4578;
  assign n4580 = A984  & ~n4563;
  assign n4581 = ~n4564 & n4580;
  assign n4582 = ~A984  & ~n4565;
  assign n4583 = ~n4581 & ~n4582;
  assign n4584 = ~n4579 & ~n4583;
  assign n4585 = ~n4575 & n4584;
  assign n4586 = ~n4574 & n4585;
  assign n4587 = ~n4574 & ~n4575;
  assign n4588 = ~n4584 & ~n4587;
  assign n4589 = ~n4586 & ~n4588;
  assign n4590 = ~n4579 & n4583;
  assign n4591 = n4579 & ~n4583;
  assign n4592 = ~n4590 & ~n4591;
  assign n4593 = n4584 & ~n4587;
  assign n4594 = ~n4567 & ~n4573;
  assign n4595 = ~n4593 & ~n4594;
  assign n4596 = ~n4592 & ~n4595;
  assign n4597 = ~n4589 & ~n4596;
  assign n4598 = ~n4589 & ~n4595;
  assign n4599 = A988  & A989 ;
  assign n4600 = A988  & ~A989 ;
  assign n4601 = ~A988  & A989 ;
  assign n4602 = ~n4600 & ~n4601;
  assign n4603 = A990  & ~n4602;
  assign n4604 = ~n4599 & ~n4603;
  assign n4605 = A985  & A986 ;
  assign n4606 = A985  & ~A986 ;
  assign n4607 = ~A985  & A986 ;
  assign n4608 = ~n4606 & ~n4607;
  assign n4609 = A987  & ~n4608;
  assign n4610 = ~n4605 & ~n4609;
  assign n4611 = ~n4604 & n4610;
  assign n4612 = n4604 & ~n4610;
  assign n4613 = ~n4611 & ~n4612;
  assign n4614 = A987  & ~n4606;
  assign n4615 = ~n4607 & n4614;
  assign n4616 = ~A987  & ~n4608;
  assign n4617 = ~n4615 & ~n4616;
  assign n4618 = A990  & ~n4600;
  assign n4619 = ~n4601 & n4618;
  assign n4620 = ~A990  & ~n4602;
  assign n4621 = ~n4619 & ~n4620;
  assign n4622 = ~n4617 & ~n4621;
  assign n4623 = ~n4613 & n4622;
  assign n4624 = ~n4604 & ~n4610;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = ~n4611 & n4622;
  assign n4627 = ~n4612 & n4626;
  assign n4628 = ~n4613 & ~n4622;
  assign n4629 = ~n4627 & ~n4628;
  assign n4630 = ~n4625 & ~n4629;
  assign n4631 = ~n4617 & n4621;
  assign n4632 = n4617 & ~n4621;
  assign n4633 = ~n4631 & ~n4632;
  assign n4634 = ~n4592 & ~n4633;
  assign n4635 = ~n4630 & n4634;
  assign n4636 = ~n4598 & n4635;
  assign n4637 = ~n4625 & ~n4633;
  assign n4638 = ~n4629 & ~n4637;
  assign n4639 = ~n4636 & ~n4638;
  assign n4640 = ~n4629 & n4634;
  assign n4641 = ~n4630 & n4640;
  assign n4642 = ~n4598 & ~n4637;
  assign n4643 = n4641 & n4642;
  assign n4644 = ~n4639 & ~n4643;
  assign n4645 = n4597 & ~n4644;
  assign n4646 = ~n4636 & n4638;
  assign n4647 = n4636 & ~n4638;
  assign n4648 = ~n4646 & ~n4647;
  assign n4649 = ~n4597 & ~n4648;
  assign n4650 = ~n4630 & ~n4633;
  assign n4651 = ~n4592 & ~n4598;
  assign n4652 = ~n4650 & n4651;
  assign n4653 = n4650 & ~n4651;
  assign n4654 = ~n4652 & ~n4653;
  assign n4655 = ~n4541 & ~n4544;
  assign n4656 = ~n4503 & ~n4509;
  assign n4657 = ~n4655 & n4656;
  assign n4658 = n4655 & ~n4656;
  assign n4659 = ~n4657 & ~n4658;
  assign n4660 = ~n4654 & ~n4659;
  assign n4661 = ~n4649 & ~n4660;
  assign n4662 = ~n4645 & n4661;
  assign n4663 = ~n4645 & ~n4649;
  assign n4664 = n4660 & ~n4663;
  assign n4665 = ~n4662 & ~n4664;
  assign n4666 = ~n4561 & ~n4665;
  assign n4667 = ~n4649 & n4660;
  assign n4668 = ~n4645 & n4667;
  assign n4669 = ~n4660 & ~n4663;
  assign n4670 = ~n4668 & ~n4669;
  assign n4671 = n4561 & ~n4670;
  assign n4672 = ~n4654 & n4659;
  assign n4673 = n4654 & ~n4659;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = ~A961  & A962 ;
  assign n4676 = A961  & ~A962 ;
  assign n4677 = A963  & ~n4676;
  assign n4678 = ~n4675 & n4677;
  assign n4679 = ~n4675 & ~n4676;
  assign n4680 = ~A963  & ~n4679;
  assign n4681 = ~n4678 & ~n4680;
  assign n4682 = ~A964  & A965 ;
  assign n4683 = A964  & ~A965 ;
  assign n4684 = A966  & ~n4683;
  assign n4685 = ~n4682 & n4684;
  assign n4686 = ~n4682 & ~n4683;
  assign n4687 = ~A966  & ~n4686;
  assign n4688 = ~n4685 & ~n4687;
  assign n4689 = ~n4681 & n4688;
  assign n4690 = n4681 & ~n4688;
  assign n4691 = ~n4689 & ~n4690;
  assign n4692 = A964  & A965 ;
  assign n4693 = A966  & ~n4686;
  assign n4694 = ~n4692 & ~n4693;
  assign n4695 = A961  & A962 ;
  assign n4696 = A963  & ~n4679;
  assign n4697 = ~n4695 & ~n4696;
  assign n4698 = ~n4694 & n4697;
  assign n4699 = n4694 & ~n4697;
  assign n4700 = ~n4698 & ~n4699;
  assign n4701 = ~n4681 & ~n4688;
  assign n4702 = ~n4700 & n4701;
  assign n4703 = ~n4694 & ~n4697;
  assign n4704 = ~n4702 & ~n4703;
  assign n4705 = ~n4698 & n4701;
  assign n4706 = ~n4699 & n4705;
  assign n4707 = ~n4700 & ~n4701;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = ~n4704 & ~n4708;
  assign n4710 = ~n4691 & ~n4709;
  assign n4711 = ~A955  & A956 ;
  assign n4712 = A955  & ~A956 ;
  assign n4713 = A957  & ~n4712;
  assign n4714 = ~n4711 & n4713;
  assign n4715 = ~n4711 & ~n4712;
  assign n4716 = ~A957  & ~n4715;
  assign n4717 = ~n4714 & ~n4716;
  assign n4718 = ~A958  & A959 ;
  assign n4719 = A958  & ~A959 ;
  assign n4720 = A960  & ~n4719;
  assign n4721 = ~n4718 & n4720;
  assign n4722 = ~n4718 & ~n4719;
  assign n4723 = ~A960  & ~n4722;
  assign n4724 = ~n4721 & ~n4723;
  assign n4725 = ~n4717 & n4724;
  assign n4726 = n4717 & ~n4724;
  assign n4727 = ~n4725 & ~n4726;
  assign n4728 = A958  & A959 ;
  assign n4729 = A960  & ~n4722;
  assign n4730 = ~n4728 & ~n4729;
  assign n4731 = A955  & A956 ;
  assign n4732 = A957  & ~n4715;
  assign n4733 = ~n4731 & ~n4732;
  assign n4734 = ~n4730 & n4733;
  assign n4735 = n4730 & ~n4733;
  assign n4736 = ~n4734 & ~n4735;
  assign n4737 = ~n4717 & ~n4724;
  assign n4738 = ~n4736 & n4737;
  assign n4739 = ~n4730 & ~n4733;
  assign n4740 = ~n4738 & ~n4739;
  assign n4741 = ~n4734 & n4737;
  assign n4742 = ~n4735 & n4741;
  assign n4743 = ~n4736 & ~n4737;
  assign n4744 = ~n4742 & ~n4743;
  assign n4745 = ~n4740 & ~n4744;
  assign n4746 = ~n4727 & ~n4745;
  assign n4747 = ~n4710 & n4746;
  assign n4748 = n4710 & ~n4746;
  assign n4749 = ~n4747 & ~n4748;
  assign n4750 = ~A949  & A950 ;
  assign n4751 = A949  & ~A950 ;
  assign n4752 = A951  & ~n4751;
  assign n4753 = ~n4750 & n4752;
  assign n4754 = ~n4750 & ~n4751;
  assign n4755 = ~A951  & ~n4754;
  assign n4756 = ~n4753 & ~n4755;
  assign n4757 = ~A952  & A953 ;
  assign n4758 = A952  & ~A953 ;
  assign n4759 = A954  & ~n4758;
  assign n4760 = ~n4757 & n4759;
  assign n4761 = ~n4757 & ~n4758;
  assign n4762 = ~A954  & ~n4761;
  assign n4763 = ~n4760 & ~n4762;
  assign n4764 = ~n4756 & n4763;
  assign n4765 = n4756 & ~n4763;
  assign n4766 = ~n4764 & ~n4765;
  assign n4767 = A952  & A953 ;
  assign n4768 = A954  & ~n4761;
  assign n4769 = ~n4767 & ~n4768;
  assign n4770 = A949  & A950 ;
  assign n4771 = A951  & ~n4754;
  assign n4772 = ~n4770 & ~n4771;
  assign n4773 = ~n4769 & n4772;
  assign n4774 = n4769 & ~n4772;
  assign n4775 = ~n4773 & ~n4774;
  assign n4776 = ~n4756 & ~n4763;
  assign n4777 = ~n4775 & n4776;
  assign n4778 = ~n4769 & ~n4772;
  assign n4779 = ~n4777 & ~n4778;
  assign n4780 = ~n4773 & n4776;
  assign n4781 = ~n4774 & n4780;
  assign n4782 = ~n4775 & ~n4776;
  assign n4783 = ~n4781 & ~n4782;
  assign n4784 = ~n4779 & ~n4783;
  assign n4785 = ~n4766 & ~n4784;
  assign n4786 = ~A943  & A944 ;
  assign n4787 = A943  & ~A944 ;
  assign n4788 = A945  & ~n4787;
  assign n4789 = ~n4786 & n4788;
  assign n4790 = ~n4786 & ~n4787;
  assign n4791 = ~A945  & ~n4790;
  assign n4792 = ~n4789 & ~n4791;
  assign n4793 = ~A946  & A947 ;
  assign n4794 = A946  & ~A947 ;
  assign n4795 = A948  & ~n4794;
  assign n4796 = ~n4793 & n4795;
  assign n4797 = ~n4793 & ~n4794;
  assign n4798 = ~A948  & ~n4797;
  assign n4799 = ~n4796 & ~n4798;
  assign n4800 = ~n4792 & n4799;
  assign n4801 = n4792 & ~n4799;
  assign n4802 = ~n4800 & ~n4801;
  assign n4803 = A946  & A947 ;
  assign n4804 = A948  & ~n4797;
  assign n4805 = ~n4803 & ~n4804;
  assign n4806 = A943  & A944 ;
  assign n4807 = A945  & ~n4790;
  assign n4808 = ~n4806 & ~n4807;
  assign n4809 = ~n4805 & n4808;
  assign n4810 = n4805 & ~n4808;
  assign n4811 = ~n4809 & ~n4810;
  assign n4812 = ~n4792 & ~n4799;
  assign n4813 = ~n4811 & n4812;
  assign n4814 = ~n4805 & ~n4808;
  assign n4815 = ~n4813 & ~n4814;
  assign n4816 = ~n4809 & n4812;
  assign n4817 = ~n4810 & n4816;
  assign n4818 = ~n4811 & ~n4812;
  assign n4819 = ~n4817 & ~n4818;
  assign n4820 = ~n4815 & ~n4819;
  assign n4821 = ~n4802 & ~n4820;
  assign n4822 = ~n4785 & n4821;
  assign n4823 = n4785 & ~n4821;
  assign n4824 = ~n4822 & ~n4823;
  assign n4825 = ~n4749 & n4824;
  assign n4826 = n4749 & ~n4824;
  assign n4827 = ~n4825 & ~n4826;
  assign n4828 = ~n4674 & ~n4827;
  assign n4829 = ~n4671 & n4828;
  assign n4830 = ~n4666 & n4829;
  assign n4831 = ~n4666 & ~n4671;
  assign n4832 = ~n4828 & ~n4831;
  assign n4833 = ~n4830 & ~n4832;
  assign n4834 = ~n4727 & ~n4740;
  assign n4835 = ~n4744 & ~n4834;
  assign n4836 = ~n4691 & ~n4727;
  assign n4837 = ~n4709 & n4836;
  assign n4838 = ~n4745 & n4837;
  assign n4839 = ~n4691 & ~n4704;
  assign n4840 = ~n4708 & ~n4839;
  assign n4841 = ~n4838 & ~n4840;
  assign n4842 = ~n4708 & n4836;
  assign n4843 = ~n4709 & n4842;
  assign n4844 = ~n4745 & ~n4839;
  assign n4845 = n4843 & n4844;
  assign n4846 = ~n4841 & ~n4845;
  assign n4847 = n4835 & ~n4846;
  assign n4848 = ~n4838 & n4840;
  assign n4849 = n4838 & ~n4840;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = ~n4835 & ~n4850;
  assign n4852 = ~n4749 & ~n4824;
  assign n4853 = ~n4851 & n4852;
  assign n4854 = ~n4847 & n4853;
  assign n4855 = ~n4847 & ~n4851;
  assign n4856 = ~n4852 & ~n4855;
  assign n4857 = ~n4854 & ~n4856;
  assign n4858 = ~n4802 & ~n4815;
  assign n4859 = ~n4819 & ~n4858;
  assign n4860 = ~n4766 & ~n4802;
  assign n4861 = ~n4784 & n4860;
  assign n4862 = ~n4820 & n4861;
  assign n4863 = ~n4766 & ~n4779;
  assign n4864 = ~n4783 & ~n4863;
  assign n4865 = ~n4862 & n4864;
  assign n4866 = n4862 & ~n4864;
  assign n4867 = ~n4865 & ~n4866;
  assign n4868 = ~n4859 & ~n4867;
  assign n4869 = ~n4862 & ~n4864;
  assign n4870 = ~n4783 & n4860;
  assign n4871 = ~n4784 & n4870;
  assign n4872 = ~n4820 & ~n4863;
  assign n4873 = n4871 & n4872;
  assign n4874 = ~n4869 & ~n4873;
  assign n4875 = n4859 & ~n4874;
  assign n4876 = ~n4868 & ~n4875;
  assign n4877 = ~n4857 & n4876;
  assign n4878 = ~n4851 & ~n4852;
  assign n4879 = ~n4847 & n4878;
  assign n4880 = n4852 & ~n4855;
  assign n4881 = ~n4879 & ~n4880;
  assign n4882 = ~n4876 & ~n4881;
  assign n4883 = ~n4877 & ~n4882;
  assign n4884 = ~n4833 & n4883;
  assign n4885 = ~n4671 & ~n4828;
  assign n4886 = ~n4666 & n4885;
  assign n4887 = n4828 & ~n4831;
  assign n4888 = ~n4886 & ~n4887;
  assign n4889 = ~n4883 & ~n4888;
  assign n4890 = ~n4884 & ~n4889;
  assign n4891 = A10  & A11 ;
  assign n4892 = A10  & ~A11 ;
  assign n4893 = ~A10  & A11 ;
  assign n4894 = ~n4892 & ~n4893;
  assign n4895 = A12  & ~n4894;
  assign n4896 = ~n4891 & ~n4895;
  assign n4897 = A7  & A8 ;
  assign n4898 = A7  & ~A8 ;
  assign n4899 = ~A7  & A8 ;
  assign n4900 = ~n4898 & ~n4899;
  assign n4901 = A9  & ~n4900;
  assign n4902 = ~n4897 & ~n4901;
  assign n4903 = n4896 & ~n4902;
  assign n4904 = ~n4896 & n4902;
  assign n4905 = A9  & ~n4898;
  assign n4906 = ~n4899 & n4905;
  assign n4907 = ~A9  & ~n4900;
  assign n4908 = ~n4906 & ~n4907;
  assign n4909 = A12  & ~n4892;
  assign n4910 = ~n4893 & n4909;
  assign n4911 = ~A12  & ~n4894;
  assign n4912 = ~n4910 & ~n4911;
  assign n4913 = ~n4908 & ~n4912;
  assign n4914 = ~n4904 & n4913;
  assign n4915 = ~n4903 & n4914;
  assign n4916 = ~n4903 & ~n4904;
  assign n4917 = ~n4913 & ~n4916;
  assign n4918 = ~n4915 & ~n4917;
  assign n4919 = ~n4908 & n4912;
  assign n4920 = n4908 & ~n4912;
  assign n4921 = ~n4919 & ~n4920;
  assign n4922 = n4913 & ~n4916;
  assign n4923 = ~n4896 & ~n4902;
  assign n4924 = ~n4922 & ~n4923;
  assign n4925 = ~n4921 & ~n4924;
  assign n4926 = ~n4918 & ~n4925;
  assign n4927 = ~n4918 & ~n4924;
  assign n4928 = A16  & A17 ;
  assign n4929 = A16  & ~A17 ;
  assign n4930 = ~A16  & A17 ;
  assign n4931 = ~n4929 & ~n4930;
  assign n4932 = A18  & ~n4931;
  assign n4933 = ~n4928 & ~n4932;
  assign n4934 = A13  & A14 ;
  assign n4935 = A13  & ~A14 ;
  assign n4936 = ~A13  & A14 ;
  assign n4937 = ~n4935 & ~n4936;
  assign n4938 = A15  & ~n4937;
  assign n4939 = ~n4934 & ~n4938;
  assign n4940 = ~n4933 & n4939;
  assign n4941 = n4933 & ~n4939;
  assign n4942 = ~n4940 & ~n4941;
  assign n4943 = A15  & ~n4935;
  assign n4944 = ~n4936 & n4943;
  assign n4945 = ~A15  & ~n4937;
  assign n4946 = ~n4944 & ~n4945;
  assign n4947 = A18  & ~n4929;
  assign n4948 = ~n4930 & n4947;
  assign n4949 = ~A18  & ~n4931;
  assign n4950 = ~n4948 & ~n4949;
  assign n4951 = ~n4946 & ~n4950;
  assign n4952 = ~n4942 & n4951;
  assign n4953 = ~n4933 & ~n4939;
  assign n4954 = ~n4952 & ~n4953;
  assign n4955 = ~n4940 & n4951;
  assign n4956 = ~n4941 & n4955;
  assign n4957 = ~n4942 & ~n4951;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = ~n4954 & ~n4958;
  assign n4960 = ~n4946 & n4950;
  assign n4961 = n4946 & ~n4950;
  assign n4962 = ~n4960 & ~n4961;
  assign n4963 = ~n4921 & ~n4962;
  assign n4964 = ~n4959 & n4963;
  assign n4965 = ~n4927 & n4964;
  assign n4966 = ~n4954 & ~n4962;
  assign n4967 = ~n4958 & ~n4966;
  assign n4968 = ~n4965 & n4967;
  assign n4969 = n4965 & ~n4967;
  assign n4970 = ~n4968 & ~n4969;
  assign n4971 = ~n4926 & ~n4970;
  assign n4972 = ~n4965 & ~n4967;
  assign n4973 = ~n4958 & n4963;
  assign n4974 = ~n4959 & n4973;
  assign n4975 = ~n4927 & ~n4966;
  assign n4976 = n4974 & n4975;
  assign n4977 = ~n4972 & ~n4976;
  assign n4978 = n4926 & ~n4977;
  assign n4979 = ~n4971 & ~n4978;
  assign n4980 = A22  & A23 ;
  assign n4981 = A22  & ~A23 ;
  assign n4982 = ~A22  & A23 ;
  assign n4983 = ~n4981 & ~n4982;
  assign n4984 = A24  & ~n4983;
  assign n4985 = ~n4980 & ~n4984;
  assign n4986 = A19  & A20 ;
  assign n4987 = A19  & ~A20 ;
  assign n4988 = ~A19  & A20 ;
  assign n4989 = ~n4987 & ~n4988;
  assign n4990 = A21  & ~n4989;
  assign n4991 = ~n4986 & ~n4990;
  assign n4992 = n4985 & ~n4991;
  assign n4993 = ~n4985 & n4991;
  assign n4994 = A21  & ~n4987;
  assign n4995 = ~n4988 & n4994;
  assign n4996 = ~A21  & ~n4989;
  assign n4997 = ~n4995 & ~n4996;
  assign n4998 = A24  & ~n4981;
  assign n4999 = ~n4982 & n4998;
  assign n5000 = ~A24  & ~n4983;
  assign n5001 = ~n4999 & ~n5000;
  assign n5002 = ~n4997 & ~n5001;
  assign n5003 = ~n4993 & n5002;
  assign n5004 = ~n4992 & n5003;
  assign n5005 = ~n4992 & ~n4993;
  assign n5006 = ~n5002 & ~n5005;
  assign n5007 = ~n5004 & ~n5006;
  assign n5008 = ~n4997 & n5001;
  assign n5009 = n4997 & ~n5001;
  assign n5010 = ~n5008 & ~n5009;
  assign n5011 = n5002 & ~n5005;
  assign n5012 = ~n4985 & ~n4991;
  assign n5013 = ~n5011 & ~n5012;
  assign n5014 = ~n5010 & ~n5013;
  assign n5015 = ~n5007 & ~n5014;
  assign n5016 = ~n5007 & ~n5013;
  assign n5017 = A28  & A29 ;
  assign n5018 = A28  & ~A29 ;
  assign n5019 = ~A28  & A29 ;
  assign n5020 = ~n5018 & ~n5019;
  assign n5021 = A30  & ~n5020;
  assign n5022 = ~n5017 & ~n5021;
  assign n5023 = A25  & A26 ;
  assign n5024 = A25  & ~A26 ;
  assign n5025 = ~A25  & A26 ;
  assign n5026 = ~n5024 & ~n5025;
  assign n5027 = A27  & ~n5026;
  assign n5028 = ~n5023 & ~n5027;
  assign n5029 = ~n5022 & n5028;
  assign n5030 = n5022 & ~n5028;
  assign n5031 = ~n5029 & ~n5030;
  assign n5032 = A27  & ~n5024;
  assign n5033 = ~n5025 & n5032;
  assign n5034 = ~A27  & ~n5026;
  assign n5035 = ~n5033 & ~n5034;
  assign n5036 = A30  & ~n5018;
  assign n5037 = ~n5019 & n5036;
  assign n5038 = ~A30  & ~n5020;
  assign n5039 = ~n5037 & ~n5038;
  assign n5040 = ~n5035 & ~n5039;
  assign n5041 = ~n5031 & n5040;
  assign n5042 = ~n5022 & ~n5028;
  assign n5043 = ~n5041 & ~n5042;
  assign n5044 = ~n5029 & n5040;
  assign n5045 = ~n5030 & n5044;
  assign n5046 = ~n5031 & ~n5040;
  assign n5047 = ~n5045 & ~n5046;
  assign n5048 = ~n5043 & ~n5047;
  assign n5049 = ~n5035 & n5039;
  assign n5050 = n5035 & ~n5039;
  assign n5051 = ~n5049 & ~n5050;
  assign n5052 = ~n5010 & ~n5051;
  assign n5053 = ~n5048 & n5052;
  assign n5054 = ~n5016 & n5053;
  assign n5055 = ~n5043 & ~n5051;
  assign n5056 = ~n5047 & ~n5055;
  assign n5057 = ~n5054 & ~n5056;
  assign n5058 = ~n5047 & n5052;
  assign n5059 = ~n5048 & n5058;
  assign n5060 = ~n5016 & ~n5055;
  assign n5061 = n5059 & n5060;
  assign n5062 = ~n5057 & ~n5061;
  assign n5063 = n5015 & ~n5062;
  assign n5064 = ~n5054 & n5056;
  assign n5065 = n5054 & ~n5056;
  assign n5066 = ~n5064 & ~n5065;
  assign n5067 = ~n5015 & ~n5066;
  assign n5068 = ~n5048 & ~n5051;
  assign n5069 = ~n5010 & ~n5016;
  assign n5070 = ~n5068 & n5069;
  assign n5071 = n5068 & ~n5069;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = ~n4959 & ~n4962;
  assign n5074 = ~n4921 & ~n4927;
  assign n5075 = ~n5073 & n5074;
  assign n5076 = n5073 & ~n5074;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = ~n5072 & ~n5077;
  assign n5079 = ~n5067 & ~n5078;
  assign n5080 = ~n5063 & n5079;
  assign n5081 = ~n5063 & ~n5067;
  assign n5082 = n5078 & ~n5081;
  assign n5083 = ~n5080 & ~n5082;
  assign n5084 = ~n4979 & ~n5083;
  assign n5085 = ~n5067 & n5078;
  assign n5086 = ~n5063 & n5085;
  assign n5087 = ~n5078 & ~n5081;
  assign n5088 = ~n5086 & ~n5087;
  assign n5089 = n4979 & ~n5088;
  assign n5090 = ~n5072 & n5077;
  assign n5091 = n5072 & ~n5077;
  assign n5092 = ~n5090 & ~n5091;
  assign n5093 = ~A991  & A992 ;
  assign n5094 = A991  & ~A992 ;
  assign n5095 = A993  & ~n5094;
  assign n5096 = ~n5093 & n5095;
  assign n5097 = ~n5093 & ~n5094;
  assign n5098 = ~A993  & ~n5097;
  assign n5099 = ~n5096 & ~n5098;
  assign n5100 = ~A994  & A995 ;
  assign n5101 = A994  & ~A995 ;
  assign n5102 = A996  & ~n5101;
  assign n5103 = ~n5100 & n5102;
  assign n5104 = ~n5100 & ~n5101;
  assign n5105 = ~A996  & ~n5104;
  assign n5106 = ~n5103 & ~n5105;
  assign n5107 = ~n5099 & n5106;
  assign n5108 = n5099 & ~n5106;
  assign n5109 = ~n5107 & ~n5108;
  assign n5110 = A994  & A995 ;
  assign n5111 = A996  & ~n5104;
  assign n5112 = ~n5110 & ~n5111;
  assign n5113 = A991  & A992 ;
  assign n5114 = A993  & ~n5097;
  assign n5115 = ~n5113 & ~n5114;
  assign n5116 = ~n5112 & n5115;
  assign n5117 = n5112 & ~n5115;
  assign n5118 = ~n5116 & ~n5117;
  assign n5119 = ~n5099 & ~n5106;
  assign n5120 = ~n5118 & n5119;
  assign n5121 = ~n5112 & ~n5115;
  assign n5122 = ~n5120 & ~n5121;
  assign n5123 = ~n5116 & n5119;
  assign n5124 = ~n5117 & n5123;
  assign n5125 = ~n5118 & ~n5119;
  assign n5126 = ~n5124 & ~n5125;
  assign n5127 = ~n5122 & ~n5126;
  assign n5128 = ~n5109 & ~n5127;
  assign n5129 = A3  & ~A4 ;
  assign n5130 = ~A3  & A4 ;
  assign n5131 = A5  & ~n5130;
  assign n5132 = ~n5129 & n5131;
  assign n5133 = ~n5129 & ~n5130;
  assign n5134 = ~A5  & ~n5133;
  assign n5135 = ~n5132 & ~n5134;
  assign n5136 = ~A0  & A1 ;
  assign n5137 = A0  & ~A1 ;
  assign n5138 = ~n5136 & ~n5137;
  assign n5139 = ~A2  & ~n5138;
  assign n5140 = A2  & ~n5136;
  assign n5141 = ~n5137 & n5140;
  assign n5142 = A6  & ~n5141;
  assign n5143 = ~n5139 & n5142;
  assign n5144 = ~n5139 & ~n5141;
  assign n5145 = ~A6  & ~n5144;
  assign n5146 = ~n5143 & ~n5145;
  assign n5147 = n5135 & ~n5146;
  assign n5148 = ~n5135 & ~n5143;
  assign n5149 = ~n5145 & n5148;
  assign n5150 = ~A997  & A998 ;
  assign n5151 = A997  & ~A998 ;
  assign n5152 = A999  & ~n5151;
  assign n5153 = ~n5150 & n5152;
  assign n5154 = ~n5150 & ~n5151;
  assign n5155 = ~A999  & ~n5154;
  assign n5156 = ~n5153 & ~n5155;
  assign n5157 = ~n5149 & ~n5156;
  assign n5158 = ~n5147 & n5157;
  assign n5159 = ~n5147 & ~n5149;
  assign n5160 = n5156 & ~n5159;
  assign n5161 = ~n5158 & ~n5160;
  assign n5162 = n5128 & n5161;
  assign n5163 = ~n5128 & ~n5161;
  assign n5164 = ~n5162 & ~n5163;
  assign n5165 = ~n5092 & ~n5164;
  assign n5166 = ~n5089 & n5165;
  assign n5167 = ~n5084 & n5166;
  assign n5168 = ~n5084 & ~n5089;
  assign n5169 = ~n5165 & ~n5168;
  assign n5170 = ~n5167 & ~n5169;
  assign n5171 = ~n5109 & ~n5122;
  assign n5172 = ~n5126 & ~n5171;
  assign n5173 = ~n5135 & ~n5146;
  assign n5174 = A6  & ~n5144;
  assign n5175 = A3  & A4 ;
  assign n5176 = A5  & ~n5133;
  assign n5177 = ~n5175 & ~n5176;
  assign n5178 = A0  & A1 ;
  assign n5179 = A2  & ~n5138;
  assign n5180 = ~n5178 & ~n5179;
  assign n5181 = ~n5177 & n5180;
  assign n5182 = n5177 & ~n5180;
  assign n5183 = ~n5181 & ~n5182;
  assign n5184 = ~n5174 & n5183;
  assign n5185 = ~n5173 & n5184;
  assign n5186 = ~n5173 & ~n5174;
  assign n5187 = ~n5183 & ~n5186;
  assign n5188 = ~n5185 & ~n5187;
  assign n5189 = ~n5156 & ~n5159;
  assign n5190 = n5188 & n5189;
  assign n5191 = A997  & A998 ;
  assign n5192 = A999  & ~n5154;
  assign n5193 = ~n5191 & ~n5192;
  assign n5194 = ~n5188 & ~n5189;
  assign n5195 = n5193 & ~n5194;
  assign n5196 = ~n5190 & n5195;
  assign n5197 = ~n5190 & ~n5194;
  assign n5198 = ~n5193 & ~n5197;
  assign n5199 = n5128 & ~n5161;
  assign n5200 = ~n5198 & n5199;
  assign n5201 = ~n5196 & n5200;
  assign n5202 = ~n5196 & ~n5198;
  assign n5203 = ~n5199 & ~n5202;
  assign n5204 = ~n5201 & ~n5203;
  assign n5205 = ~n5172 & ~n5204;
  assign n5206 = ~n5198 & ~n5199;
  assign n5207 = ~n5196 & n5206;
  assign n5208 = n5199 & ~n5202;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = n5172 & ~n5209;
  assign n5211 = ~n5205 & ~n5210;
  assign n5212 = ~n5170 & n5211;
  assign n5213 = ~n5089 & ~n5165;
  assign n5214 = ~n5084 & n5213;
  assign n5215 = n5165 & ~n5168;
  assign n5216 = ~n5214 & ~n5215;
  assign n5217 = ~n5211 & ~n5216;
  assign n5218 = ~n5212 & ~n5217;
  assign n5219 = A46  & A47 ;
  assign n5220 = A46  & ~A47 ;
  assign n5221 = ~A46  & A47 ;
  assign n5222 = ~n5220 & ~n5221;
  assign n5223 = A48  & ~n5222;
  assign n5224 = ~n5219 & ~n5223;
  assign n5225 = A43  & A44 ;
  assign n5226 = A43  & ~A44 ;
  assign n5227 = ~A43  & A44 ;
  assign n5228 = ~n5226 & ~n5227;
  assign n5229 = A45  & ~n5228;
  assign n5230 = ~n5225 & ~n5229;
  assign n5231 = n5224 & ~n5230;
  assign n5232 = ~n5224 & n5230;
  assign n5233 = A45  & ~n5226;
  assign n5234 = ~n5227 & n5233;
  assign n5235 = ~A45  & ~n5228;
  assign n5236 = ~n5234 & ~n5235;
  assign n5237 = A48  & ~n5220;
  assign n5238 = ~n5221 & n5237;
  assign n5239 = ~A48  & ~n5222;
  assign n5240 = ~n5238 & ~n5239;
  assign n5241 = ~n5236 & ~n5240;
  assign n5242 = ~n5232 & n5241;
  assign n5243 = ~n5231 & n5242;
  assign n5244 = ~n5231 & ~n5232;
  assign n5245 = ~n5241 & ~n5244;
  assign n5246 = ~n5243 & ~n5245;
  assign n5247 = ~n5236 & n5240;
  assign n5248 = n5236 & ~n5240;
  assign n5249 = ~n5247 & ~n5248;
  assign n5250 = n5241 & ~n5244;
  assign n5251 = ~n5224 & ~n5230;
  assign n5252 = ~n5250 & ~n5251;
  assign n5253 = ~n5249 & ~n5252;
  assign n5254 = ~n5246 & ~n5253;
  assign n5255 = ~n5246 & ~n5252;
  assign n5256 = A52  & A53 ;
  assign n5257 = A52  & ~A53 ;
  assign n5258 = ~A52  & A53 ;
  assign n5259 = ~n5257 & ~n5258;
  assign n5260 = A54  & ~n5259;
  assign n5261 = ~n5256 & ~n5260;
  assign n5262 = A49  & A50 ;
  assign n5263 = A49  & ~A50 ;
  assign n5264 = ~A49  & A50 ;
  assign n5265 = ~n5263 & ~n5264;
  assign n5266 = A51  & ~n5265;
  assign n5267 = ~n5262 & ~n5266;
  assign n5268 = ~n5261 & n5267;
  assign n5269 = n5261 & ~n5267;
  assign n5270 = ~n5268 & ~n5269;
  assign n5271 = A51  & ~n5263;
  assign n5272 = ~n5264 & n5271;
  assign n5273 = ~A51  & ~n5265;
  assign n5274 = ~n5272 & ~n5273;
  assign n5275 = A54  & ~n5257;
  assign n5276 = ~n5258 & n5275;
  assign n5277 = ~A54  & ~n5259;
  assign n5278 = ~n5276 & ~n5277;
  assign n5279 = ~n5274 & ~n5278;
  assign n5280 = ~n5270 & n5279;
  assign n5281 = ~n5261 & ~n5267;
  assign n5282 = ~n5280 & ~n5281;
  assign n5283 = ~n5268 & n5279;
  assign n5284 = ~n5269 & n5283;
  assign n5285 = ~n5270 & ~n5279;
  assign n5286 = ~n5284 & ~n5285;
  assign n5287 = ~n5282 & ~n5286;
  assign n5288 = ~n5274 & n5278;
  assign n5289 = n5274 & ~n5278;
  assign n5290 = ~n5288 & ~n5289;
  assign n5291 = ~n5249 & ~n5290;
  assign n5292 = ~n5287 & n5291;
  assign n5293 = ~n5255 & n5292;
  assign n5294 = ~n5282 & ~n5290;
  assign n5295 = ~n5286 & ~n5294;
  assign n5296 = ~n5293 & ~n5295;
  assign n5297 = ~n5286 & n5291;
  assign n5298 = ~n5287 & n5297;
  assign n5299 = ~n5255 & ~n5294;
  assign n5300 = n5298 & n5299;
  assign n5301 = ~n5296 & ~n5300;
  assign n5302 = n5254 & ~n5301;
  assign n5303 = ~n5293 & n5295;
  assign n5304 = n5293 & ~n5295;
  assign n5305 = ~n5303 & ~n5304;
  assign n5306 = ~n5254 & ~n5305;
  assign n5307 = ~n5287 & ~n5290;
  assign n5308 = ~n5249 & ~n5255;
  assign n5309 = ~n5307 & n5308;
  assign n5310 = n5307 & ~n5308;
  assign n5311 = ~n5309 & ~n5310;
  assign n5312 = ~A37  & A38 ;
  assign n5313 = A37  & ~A38 ;
  assign n5314 = A39  & ~n5313;
  assign n5315 = ~n5312 & n5314;
  assign n5316 = ~n5312 & ~n5313;
  assign n5317 = ~A39  & ~n5316;
  assign n5318 = ~n5315 & ~n5317;
  assign n5319 = ~A40  & A41 ;
  assign n5320 = A40  & ~A41 ;
  assign n5321 = A42  & ~n5320;
  assign n5322 = ~n5319 & n5321;
  assign n5323 = ~n5319 & ~n5320;
  assign n5324 = ~A42  & ~n5323;
  assign n5325 = ~n5322 & ~n5324;
  assign n5326 = ~n5318 & n5325;
  assign n5327 = n5318 & ~n5325;
  assign n5328 = ~n5326 & ~n5327;
  assign n5329 = A40  & A41 ;
  assign n5330 = A42  & ~n5323;
  assign n5331 = ~n5329 & ~n5330;
  assign n5332 = A37  & A38 ;
  assign n5333 = A39  & ~n5316;
  assign n5334 = ~n5332 & ~n5333;
  assign n5335 = ~n5331 & n5334;
  assign n5336 = n5331 & ~n5334;
  assign n5337 = ~n5335 & ~n5336;
  assign n5338 = ~n5318 & ~n5325;
  assign n5339 = ~n5337 & n5338;
  assign n5340 = ~n5331 & ~n5334;
  assign n5341 = ~n5339 & ~n5340;
  assign n5342 = ~n5335 & n5338;
  assign n5343 = ~n5336 & n5342;
  assign n5344 = ~n5337 & ~n5338;
  assign n5345 = ~n5343 & ~n5344;
  assign n5346 = ~n5341 & ~n5345;
  assign n5347 = ~n5328 & ~n5346;
  assign n5348 = ~A31  & A32 ;
  assign n5349 = A31  & ~A32 ;
  assign n5350 = A33  & ~n5349;
  assign n5351 = ~n5348 & n5350;
  assign n5352 = ~n5348 & ~n5349;
  assign n5353 = ~A33  & ~n5352;
  assign n5354 = ~n5351 & ~n5353;
  assign n5355 = ~A34  & A35 ;
  assign n5356 = A34  & ~A35 ;
  assign n5357 = A36  & ~n5356;
  assign n5358 = ~n5355 & n5357;
  assign n5359 = ~n5355 & ~n5356;
  assign n5360 = ~A36  & ~n5359;
  assign n5361 = ~n5358 & ~n5360;
  assign n5362 = ~n5354 & n5361;
  assign n5363 = n5354 & ~n5361;
  assign n5364 = ~n5362 & ~n5363;
  assign n5365 = A34  & A35 ;
  assign n5366 = A36  & ~n5359;
  assign n5367 = ~n5365 & ~n5366;
  assign n5368 = A31  & A32 ;
  assign n5369 = A33  & ~n5352;
  assign n5370 = ~n5368 & ~n5369;
  assign n5371 = ~n5367 & n5370;
  assign n5372 = n5367 & ~n5370;
  assign n5373 = ~n5371 & ~n5372;
  assign n5374 = ~n5354 & ~n5361;
  assign n5375 = ~n5373 & n5374;
  assign n5376 = ~n5367 & ~n5370;
  assign n5377 = ~n5375 & ~n5376;
  assign n5378 = ~n5371 & n5374;
  assign n5379 = ~n5372 & n5378;
  assign n5380 = ~n5373 & ~n5374;
  assign n5381 = ~n5379 & ~n5380;
  assign n5382 = ~n5377 & ~n5381;
  assign n5383 = ~n5364 & ~n5382;
  assign n5384 = ~n5347 & n5383;
  assign n5385 = n5347 & ~n5383;
  assign n5386 = ~n5384 & ~n5385;
  assign n5387 = ~n5311 & ~n5386;
  assign n5388 = ~n5306 & n5387;
  assign n5389 = ~n5302 & n5388;
  assign n5390 = ~n5302 & ~n5306;
  assign n5391 = ~n5387 & ~n5390;
  assign n5392 = ~n5389 & ~n5391;
  assign n5393 = ~n5364 & ~n5377;
  assign n5394 = ~n5381 & ~n5393;
  assign n5395 = ~n5328 & ~n5364;
  assign n5396 = ~n5346 & n5395;
  assign n5397 = ~n5382 & n5396;
  assign n5398 = ~n5328 & ~n5341;
  assign n5399 = ~n5345 & ~n5398;
  assign n5400 = ~n5397 & n5399;
  assign n5401 = n5397 & ~n5399;
  assign n5402 = ~n5400 & ~n5401;
  assign n5403 = ~n5394 & ~n5402;
  assign n5404 = ~n5397 & ~n5399;
  assign n5405 = ~n5345 & n5395;
  assign n5406 = ~n5346 & n5405;
  assign n5407 = ~n5382 & ~n5398;
  assign n5408 = n5406 & n5407;
  assign n5409 = ~n5404 & ~n5408;
  assign n5410 = n5394 & ~n5409;
  assign n5411 = ~n5403 & ~n5410;
  assign n5412 = ~n5392 & n5411;
  assign n5413 = ~n5306 & ~n5387;
  assign n5414 = ~n5302 & n5413;
  assign n5415 = n5387 & ~n5390;
  assign n5416 = ~n5414 & ~n5415;
  assign n5417 = ~n5411 & ~n5416;
  assign n5418 = ~n5412 & ~n5417;
  assign n5419 = A58  & A59 ;
  assign n5420 = A58  & ~A59 ;
  assign n5421 = ~A58  & A59 ;
  assign n5422 = ~n5420 & ~n5421;
  assign n5423 = A60  & ~n5422;
  assign n5424 = ~n5419 & ~n5423;
  assign n5425 = A55  & A56 ;
  assign n5426 = A55  & ~A56 ;
  assign n5427 = ~A55  & A56 ;
  assign n5428 = ~n5426 & ~n5427;
  assign n5429 = A57  & ~n5428;
  assign n5430 = ~n5425 & ~n5429;
  assign n5431 = n5424 & ~n5430;
  assign n5432 = ~n5424 & n5430;
  assign n5433 = A57  & ~n5426;
  assign n5434 = ~n5427 & n5433;
  assign n5435 = ~A57  & ~n5428;
  assign n5436 = ~n5434 & ~n5435;
  assign n5437 = A60  & ~n5420;
  assign n5438 = ~n5421 & n5437;
  assign n5439 = ~A60  & ~n5422;
  assign n5440 = ~n5438 & ~n5439;
  assign n5441 = ~n5436 & ~n5440;
  assign n5442 = ~n5432 & n5441;
  assign n5443 = ~n5431 & n5442;
  assign n5444 = ~n5431 & ~n5432;
  assign n5445 = ~n5441 & ~n5444;
  assign n5446 = ~n5443 & ~n5445;
  assign n5447 = ~n5436 & n5440;
  assign n5448 = n5436 & ~n5440;
  assign n5449 = ~n5447 & ~n5448;
  assign n5450 = n5441 & ~n5444;
  assign n5451 = ~n5424 & ~n5430;
  assign n5452 = ~n5450 & ~n5451;
  assign n5453 = ~n5449 & ~n5452;
  assign n5454 = ~n5446 & ~n5453;
  assign n5455 = ~n5446 & ~n5452;
  assign n5456 = A64  & A65 ;
  assign n5457 = A64  & ~A65 ;
  assign n5458 = ~A64  & A65 ;
  assign n5459 = ~n5457 & ~n5458;
  assign n5460 = A66  & ~n5459;
  assign n5461 = ~n5456 & ~n5460;
  assign n5462 = A61  & A62 ;
  assign n5463 = A61  & ~A62 ;
  assign n5464 = ~A61  & A62 ;
  assign n5465 = ~n5463 & ~n5464;
  assign n5466 = A63  & ~n5465;
  assign n5467 = ~n5462 & ~n5466;
  assign n5468 = ~n5461 & n5467;
  assign n5469 = n5461 & ~n5467;
  assign n5470 = ~n5468 & ~n5469;
  assign n5471 = A63  & ~n5463;
  assign n5472 = ~n5464 & n5471;
  assign n5473 = ~A63  & ~n5465;
  assign n5474 = ~n5472 & ~n5473;
  assign n5475 = A66  & ~n5457;
  assign n5476 = ~n5458 & n5475;
  assign n5477 = ~A66  & ~n5459;
  assign n5478 = ~n5476 & ~n5477;
  assign n5479 = ~n5474 & ~n5478;
  assign n5480 = ~n5470 & n5479;
  assign n5481 = ~n5461 & ~n5467;
  assign n5482 = ~n5480 & ~n5481;
  assign n5483 = ~n5468 & n5479;
  assign n5484 = ~n5469 & n5483;
  assign n5485 = ~n5470 & ~n5479;
  assign n5486 = ~n5484 & ~n5485;
  assign n5487 = ~n5482 & ~n5486;
  assign n5488 = ~n5474 & n5478;
  assign n5489 = n5474 & ~n5478;
  assign n5490 = ~n5488 & ~n5489;
  assign n5491 = ~n5449 & ~n5490;
  assign n5492 = ~n5487 & n5491;
  assign n5493 = ~n5455 & n5492;
  assign n5494 = ~n5482 & ~n5490;
  assign n5495 = ~n5486 & ~n5494;
  assign n5496 = ~n5493 & n5495;
  assign n5497 = n5493 & ~n5495;
  assign n5498 = ~n5496 & ~n5497;
  assign n5499 = ~n5454 & ~n5498;
  assign n5500 = ~n5493 & ~n5495;
  assign n5501 = ~n5486 & n5491;
  assign n5502 = ~n5487 & n5501;
  assign n5503 = ~n5455 & ~n5494;
  assign n5504 = n5502 & n5503;
  assign n5505 = ~n5500 & ~n5504;
  assign n5506 = n5454 & ~n5505;
  assign n5507 = ~n5499 & ~n5506;
  assign n5508 = A70  & A71 ;
  assign n5509 = A70  & ~A71 ;
  assign n5510 = ~A70  & A71 ;
  assign n5511 = ~n5509 & ~n5510;
  assign n5512 = A72  & ~n5511;
  assign n5513 = ~n5508 & ~n5512;
  assign n5514 = A67  & A68 ;
  assign n5515 = A67  & ~A68 ;
  assign n5516 = ~A67  & A68 ;
  assign n5517 = ~n5515 & ~n5516;
  assign n5518 = A69  & ~n5517;
  assign n5519 = ~n5514 & ~n5518;
  assign n5520 = n5513 & ~n5519;
  assign n5521 = ~n5513 & n5519;
  assign n5522 = A69  & ~n5515;
  assign n5523 = ~n5516 & n5522;
  assign n5524 = ~A69  & ~n5517;
  assign n5525 = ~n5523 & ~n5524;
  assign n5526 = A72  & ~n5509;
  assign n5527 = ~n5510 & n5526;
  assign n5528 = ~A72  & ~n5511;
  assign n5529 = ~n5527 & ~n5528;
  assign n5530 = ~n5525 & ~n5529;
  assign n5531 = ~n5521 & n5530;
  assign n5532 = ~n5520 & n5531;
  assign n5533 = ~n5520 & ~n5521;
  assign n5534 = ~n5530 & ~n5533;
  assign n5535 = ~n5532 & ~n5534;
  assign n5536 = ~n5525 & n5529;
  assign n5537 = n5525 & ~n5529;
  assign n5538 = ~n5536 & ~n5537;
  assign n5539 = n5530 & ~n5533;
  assign n5540 = ~n5513 & ~n5519;
  assign n5541 = ~n5539 & ~n5540;
  assign n5542 = ~n5538 & ~n5541;
  assign n5543 = ~n5535 & ~n5542;
  assign n5544 = ~n5535 & ~n5541;
  assign n5545 = A76  & A77 ;
  assign n5546 = A76  & ~A77 ;
  assign n5547 = ~A76  & A77 ;
  assign n5548 = ~n5546 & ~n5547;
  assign n5549 = A78  & ~n5548;
  assign n5550 = ~n5545 & ~n5549;
  assign n5551 = A73  & A74 ;
  assign n5552 = A73  & ~A74 ;
  assign n5553 = ~A73  & A74 ;
  assign n5554 = ~n5552 & ~n5553;
  assign n5555 = A75  & ~n5554;
  assign n5556 = ~n5551 & ~n5555;
  assign n5557 = ~n5550 & n5556;
  assign n5558 = n5550 & ~n5556;
  assign n5559 = ~n5557 & ~n5558;
  assign n5560 = A75  & ~n5552;
  assign n5561 = ~n5553 & n5560;
  assign n5562 = ~A75  & ~n5554;
  assign n5563 = ~n5561 & ~n5562;
  assign n5564 = A78  & ~n5546;
  assign n5565 = ~n5547 & n5564;
  assign n5566 = ~A78  & ~n5548;
  assign n5567 = ~n5565 & ~n5566;
  assign n5568 = ~n5563 & ~n5567;
  assign n5569 = ~n5559 & n5568;
  assign n5570 = ~n5550 & ~n5556;
  assign n5571 = ~n5569 & ~n5570;
  assign n5572 = ~n5557 & n5568;
  assign n5573 = ~n5558 & n5572;
  assign n5574 = ~n5559 & ~n5568;
  assign n5575 = ~n5573 & ~n5574;
  assign n5576 = ~n5571 & ~n5575;
  assign n5577 = ~n5563 & n5567;
  assign n5578 = n5563 & ~n5567;
  assign n5579 = ~n5577 & ~n5578;
  assign n5580 = ~n5538 & ~n5579;
  assign n5581 = ~n5576 & n5580;
  assign n5582 = ~n5544 & n5581;
  assign n5583 = ~n5571 & ~n5579;
  assign n5584 = ~n5575 & ~n5583;
  assign n5585 = ~n5582 & ~n5584;
  assign n5586 = ~n5575 & n5580;
  assign n5587 = ~n5576 & n5586;
  assign n5588 = ~n5544 & ~n5583;
  assign n5589 = n5587 & n5588;
  assign n5590 = ~n5585 & ~n5589;
  assign n5591 = n5543 & ~n5590;
  assign n5592 = ~n5582 & n5584;
  assign n5593 = n5582 & ~n5584;
  assign n5594 = ~n5592 & ~n5593;
  assign n5595 = ~n5543 & ~n5594;
  assign n5596 = ~n5576 & ~n5579;
  assign n5597 = ~n5538 & ~n5544;
  assign n5598 = ~n5596 & n5597;
  assign n5599 = n5596 & ~n5597;
  assign n5600 = ~n5598 & ~n5599;
  assign n5601 = ~n5487 & ~n5490;
  assign n5602 = ~n5449 & ~n5455;
  assign n5603 = ~n5601 & n5602;
  assign n5604 = n5601 & ~n5602;
  assign n5605 = ~n5603 & ~n5604;
  assign n5606 = ~n5600 & ~n5605;
  assign n5607 = ~n5595 & ~n5606;
  assign n5608 = ~n5591 & n5607;
  assign n5609 = ~n5591 & ~n5595;
  assign n5610 = n5606 & ~n5609;
  assign n5611 = ~n5608 & ~n5610;
  assign n5612 = ~n5507 & ~n5611;
  assign n5613 = ~n5595 & n5606;
  assign n5614 = ~n5591 & n5613;
  assign n5615 = ~n5606 & ~n5609;
  assign n5616 = ~n5614 & ~n5615;
  assign n5617 = n5507 & ~n5616;
  assign n5618 = ~n5600 & n5605;
  assign n5619 = n5600 & ~n5605;
  assign n5620 = ~n5618 & ~n5619;
  assign n5621 = ~n5311 & n5386;
  assign n5622 = n5311 & ~n5386;
  assign n5623 = ~n5621 & ~n5622;
  assign n5624 = ~n5620 & ~n5623;
  assign n5625 = ~n5617 & ~n5624;
  assign n5626 = ~n5612 & n5625;
  assign n5627 = ~n5612 & ~n5617;
  assign n5628 = n5624 & ~n5627;
  assign n5629 = ~n5626 & ~n5628;
  assign n5630 = ~n5418 & ~n5629;
  assign n5631 = ~n5617 & n5624;
  assign n5632 = ~n5612 & n5631;
  assign n5633 = ~n5624 & ~n5627;
  assign n5634 = ~n5632 & ~n5633;
  assign n5635 = n5418 & ~n5634;
  assign n5636 = ~n5620 & n5623;
  assign n5637 = n5620 & ~n5623;
  assign n5638 = ~n5636 & ~n5637;
  assign n5639 = ~n5092 & n5164;
  assign n5640 = ~n5090 & ~n5164;
  assign n5641 = ~n5091 & n5640;
  assign n5642 = ~n5639 & ~n5641;
  assign n5643 = ~n5638 & ~n5642;
  assign n5644 = ~n5635 & ~n5643;
  assign n5645 = ~n5630 & n5644;
  assign n5646 = ~n5630 & ~n5635;
  assign n5647 = n5643 & ~n5646;
  assign n5648 = ~n5645 & ~n5647;
  assign n5649 = ~n5218 & ~n5648;
  assign n5650 = ~n5635 & n5643;
  assign n5651 = ~n5630 & n5650;
  assign n5652 = ~n5643 & ~n5646;
  assign n5653 = ~n5651 & ~n5652;
  assign n5654 = n5218 & ~n5653;
  assign n5655 = ~n5638 & n5642;
  assign n5656 = n5638 & ~n5642;
  assign n5657 = ~n5655 & ~n5656;
  assign n5658 = ~n4674 & n4827;
  assign n5659 = n4674 & ~n4827;
  assign n5660 = ~n5658 & ~n5659;
  assign n5661 = ~n5657 & ~n5660;
  assign n5662 = ~n5654 & ~n5661;
  assign n5663 = ~n5649 & n5662;
  assign n5664 = ~n5649 & ~n5654;
  assign n5665 = n5661 & ~n5664;
  assign n5666 = ~n5663 & ~n5665;
  assign n5667 = ~n4890 & ~n5666;
  assign n5668 = ~n5654 & n5661;
  assign n5669 = ~n5649 & n5668;
  assign n5670 = ~n5661 & ~n5664;
  assign n5671 = ~n5669 & ~n5670;
  assign n5672 = n4890 & ~n5671;
  assign n5673 = ~n5657 & n5660;
  assign n5674 = ~n5655 & ~n5660;
  assign n5675 = ~n5656 & n5674;
  assign n5676 = ~n5673 & ~n5675;
  assign n5677 = ~A937  & A938 ;
  assign n5678 = A937  & ~A938 ;
  assign n5679 = A939  & ~n5678;
  assign n5680 = ~n5677 & n5679;
  assign n5681 = ~n5677 & ~n5678;
  assign n5682 = ~A939  & ~n5681;
  assign n5683 = ~n5680 & ~n5682;
  assign n5684 = ~A940  & A941 ;
  assign n5685 = A940  & ~A941 ;
  assign n5686 = A942  & ~n5685;
  assign n5687 = ~n5684 & n5686;
  assign n5688 = ~n5684 & ~n5685;
  assign n5689 = ~A942  & ~n5688;
  assign n5690 = ~n5687 & ~n5689;
  assign n5691 = ~n5683 & n5690;
  assign n5692 = n5683 & ~n5690;
  assign n5693 = ~n5691 & ~n5692;
  assign n5694 = A940  & A941 ;
  assign n5695 = A942  & ~n5688;
  assign n5696 = ~n5694 & ~n5695;
  assign n5697 = A937  & A938 ;
  assign n5698 = A939  & ~n5681;
  assign n5699 = ~n5697 & ~n5698;
  assign n5700 = ~n5696 & n5699;
  assign n5701 = n5696 & ~n5699;
  assign n5702 = ~n5700 & ~n5701;
  assign n5703 = ~n5683 & ~n5690;
  assign n5704 = ~n5702 & n5703;
  assign n5705 = ~n5696 & ~n5699;
  assign n5706 = ~n5704 & ~n5705;
  assign n5707 = ~n5700 & n5703;
  assign n5708 = ~n5701 & n5707;
  assign n5709 = ~n5702 & ~n5703;
  assign n5710 = ~n5708 & ~n5709;
  assign n5711 = ~n5706 & ~n5710;
  assign n5712 = ~n5693 & ~n5711;
  assign n5713 = ~A931  & A932 ;
  assign n5714 = A931  & ~A932 ;
  assign n5715 = A933  & ~n5714;
  assign n5716 = ~n5713 & n5715;
  assign n5717 = ~n5713 & ~n5714;
  assign n5718 = ~A933  & ~n5717;
  assign n5719 = ~n5716 & ~n5718;
  assign n5720 = ~A934  & A935 ;
  assign n5721 = A934  & ~A935 ;
  assign n5722 = A936  & ~n5721;
  assign n5723 = ~n5720 & n5722;
  assign n5724 = ~n5720 & ~n5721;
  assign n5725 = ~A936  & ~n5724;
  assign n5726 = ~n5723 & ~n5725;
  assign n5727 = ~n5719 & n5726;
  assign n5728 = n5719 & ~n5726;
  assign n5729 = ~n5727 & ~n5728;
  assign n5730 = A934  & A935 ;
  assign n5731 = A936  & ~n5724;
  assign n5732 = ~n5730 & ~n5731;
  assign n5733 = A931  & A932 ;
  assign n5734 = A933  & ~n5717;
  assign n5735 = ~n5733 & ~n5734;
  assign n5736 = ~n5732 & n5735;
  assign n5737 = n5732 & ~n5735;
  assign n5738 = ~n5736 & ~n5737;
  assign n5739 = ~n5719 & ~n5726;
  assign n5740 = ~n5738 & n5739;
  assign n5741 = ~n5732 & ~n5735;
  assign n5742 = ~n5740 & ~n5741;
  assign n5743 = ~n5736 & n5739;
  assign n5744 = ~n5737 & n5743;
  assign n5745 = ~n5738 & ~n5739;
  assign n5746 = ~n5744 & ~n5745;
  assign n5747 = ~n5742 & ~n5746;
  assign n5748 = ~n5729 & ~n5747;
  assign n5749 = ~n5712 & n5748;
  assign n5750 = n5712 & ~n5748;
  assign n5751 = ~n5749 & ~n5750;
  assign n5752 = ~A925  & A926 ;
  assign n5753 = A925  & ~A926 ;
  assign n5754 = A927  & ~n5753;
  assign n5755 = ~n5752 & n5754;
  assign n5756 = ~n5752 & ~n5753;
  assign n5757 = ~A927  & ~n5756;
  assign n5758 = ~n5755 & ~n5757;
  assign n5759 = ~A928  & A929 ;
  assign n5760 = A928  & ~A929 ;
  assign n5761 = A930  & ~n5760;
  assign n5762 = ~n5759 & n5761;
  assign n5763 = ~n5759 & ~n5760;
  assign n5764 = ~A930  & ~n5763;
  assign n5765 = ~n5762 & ~n5764;
  assign n5766 = ~n5758 & n5765;
  assign n5767 = n5758 & ~n5765;
  assign n5768 = ~n5766 & ~n5767;
  assign n5769 = A928  & A929 ;
  assign n5770 = A930  & ~n5763;
  assign n5771 = ~n5769 & ~n5770;
  assign n5772 = A925  & A926 ;
  assign n5773 = A927  & ~n5756;
  assign n5774 = ~n5772 & ~n5773;
  assign n5775 = ~n5771 & n5774;
  assign n5776 = n5771 & ~n5774;
  assign n5777 = ~n5775 & ~n5776;
  assign n5778 = ~n5758 & ~n5765;
  assign n5779 = ~n5777 & n5778;
  assign n5780 = ~n5771 & ~n5774;
  assign n5781 = ~n5779 & ~n5780;
  assign n5782 = ~n5775 & n5778;
  assign n5783 = ~n5776 & n5782;
  assign n5784 = ~n5777 & ~n5778;
  assign n5785 = ~n5783 & ~n5784;
  assign n5786 = ~n5781 & ~n5785;
  assign n5787 = ~n5768 & ~n5786;
  assign n5788 = ~A919  & A920 ;
  assign n5789 = A919  & ~A920 ;
  assign n5790 = A921  & ~n5789;
  assign n5791 = ~n5788 & n5790;
  assign n5792 = ~n5788 & ~n5789;
  assign n5793 = ~A921  & ~n5792;
  assign n5794 = ~n5791 & ~n5793;
  assign n5795 = ~A922  & A923 ;
  assign n5796 = A922  & ~A923 ;
  assign n5797 = A924  & ~n5796;
  assign n5798 = ~n5795 & n5797;
  assign n5799 = ~n5795 & ~n5796;
  assign n5800 = ~A924  & ~n5799;
  assign n5801 = ~n5798 & ~n5800;
  assign n5802 = ~n5794 & n5801;
  assign n5803 = n5794 & ~n5801;
  assign n5804 = ~n5802 & ~n5803;
  assign n5805 = A922  & A923 ;
  assign n5806 = A924  & ~n5799;
  assign n5807 = ~n5805 & ~n5806;
  assign n5808 = A919  & A920 ;
  assign n5809 = A921  & ~n5792;
  assign n5810 = ~n5808 & ~n5809;
  assign n5811 = ~n5807 & n5810;
  assign n5812 = n5807 & ~n5810;
  assign n5813 = ~n5811 & ~n5812;
  assign n5814 = ~n5794 & ~n5801;
  assign n5815 = ~n5813 & n5814;
  assign n5816 = ~n5807 & ~n5810;
  assign n5817 = ~n5815 & ~n5816;
  assign n5818 = ~n5811 & n5814;
  assign n5819 = ~n5812 & n5818;
  assign n5820 = ~n5813 & ~n5814;
  assign n5821 = ~n5819 & ~n5820;
  assign n5822 = ~n5817 & ~n5821;
  assign n5823 = ~n5804 & ~n5822;
  assign n5824 = ~n5787 & n5823;
  assign n5825 = n5787 & ~n5823;
  assign n5826 = ~n5824 & ~n5825;
  assign n5827 = ~n5751 & n5826;
  assign n5828 = n5751 & ~n5826;
  assign n5829 = ~n5827 & ~n5828;
  assign n5830 = ~A913  & A914 ;
  assign n5831 = A913  & ~A914 ;
  assign n5832 = A915  & ~n5831;
  assign n5833 = ~n5830 & n5832;
  assign n5834 = ~n5830 & ~n5831;
  assign n5835 = ~A915  & ~n5834;
  assign n5836 = ~n5833 & ~n5835;
  assign n5837 = ~A916  & A917 ;
  assign n5838 = A916  & ~A917 ;
  assign n5839 = A918  & ~n5838;
  assign n5840 = ~n5837 & n5839;
  assign n5841 = ~n5837 & ~n5838;
  assign n5842 = ~A918  & ~n5841;
  assign n5843 = ~n5840 & ~n5842;
  assign n5844 = ~n5836 & n5843;
  assign n5845 = n5836 & ~n5843;
  assign n5846 = ~n5844 & ~n5845;
  assign n5847 = A916  & A917 ;
  assign n5848 = A918  & ~n5841;
  assign n5849 = ~n5847 & ~n5848;
  assign n5850 = A913  & A914 ;
  assign n5851 = A915  & ~n5834;
  assign n5852 = ~n5850 & ~n5851;
  assign n5853 = ~n5849 & n5852;
  assign n5854 = n5849 & ~n5852;
  assign n5855 = ~n5853 & ~n5854;
  assign n5856 = ~n5836 & ~n5843;
  assign n5857 = ~n5855 & n5856;
  assign n5858 = ~n5849 & ~n5852;
  assign n5859 = ~n5857 & ~n5858;
  assign n5860 = ~n5853 & n5856;
  assign n5861 = ~n5854 & n5860;
  assign n5862 = ~n5855 & ~n5856;
  assign n5863 = ~n5861 & ~n5862;
  assign n5864 = ~n5859 & ~n5863;
  assign n5865 = ~n5846 & ~n5864;
  assign n5866 = ~A907  & A908 ;
  assign n5867 = A907  & ~A908 ;
  assign n5868 = A909  & ~n5867;
  assign n5869 = ~n5866 & n5868;
  assign n5870 = ~n5866 & ~n5867;
  assign n5871 = ~A909  & ~n5870;
  assign n5872 = ~n5869 & ~n5871;
  assign n5873 = ~A910  & A911 ;
  assign n5874 = A910  & ~A911 ;
  assign n5875 = A912  & ~n5874;
  assign n5876 = ~n5873 & n5875;
  assign n5877 = ~n5873 & ~n5874;
  assign n5878 = ~A912  & ~n5877;
  assign n5879 = ~n5876 & ~n5878;
  assign n5880 = ~n5872 & n5879;
  assign n5881 = n5872 & ~n5879;
  assign n5882 = ~n5880 & ~n5881;
  assign n5883 = A910  & A911 ;
  assign n5884 = A912  & ~n5877;
  assign n5885 = ~n5883 & ~n5884;
  assign n5886 = A907  & A908 ;
  assign n5887 = A909  & ~n5870;
  assign n5888 = ~n5886 & ~n5887;
  assign n5889 = ~n5885 & n5888;
  assign n5890 = n5885 & ~n5888;
  assign n5891 = ~n5889 & ~n5890;
  assign n5892 = ~n5872 & ~n5879;
  assign n5893 = ~n5891 & n5892;
  assign n5894 = ~n5885 & ~n5888;
  assign n5895 = ~n5893 & ~n5894;
  assign n5896 = ~n5889 & n5892;
  assign n5897 = ~n5890 & n5896;
  assign n5898 = ~n5891 & ~n5892;
  assign n5899 = ~n5897 & ~n5898;
  assign n5900 = ~n5895 & ~n5899;
  assign n5901 = ~n5882 & ~n5900;
  assign n5902 = ~n5865 & n5901;
  assign n5903 = n5865 & ~n5901;
  assign n5904 = ~n5902 & ~n5903;
  assign n5905 = ~A901  & A902 ;
  assign n5906 = A901  & ~A902 ;
  assign n5907 = A903  & ~n5906;
  assign n5908 = ~n5905 & n5907;
  assign n5909 = ~n5905 & ~n5906;
  assign n5910 = ~A903  & ~n5909;
  assign n5911 = ~n5908 & ~n5910;
  assign n5912 = ~A904  & A905 ;
  assign n5913 = A904  & ~A905 ;
  assign n5914 = A906  & ~n5913;
  assign n5915 = ~n5912 & n5914;
  assign n5916 = ~n5912 & ~n5913;
  assign n5917 = ~A906  & ~n5916;
  assign n5918 = ~n5915 & ~n5917;
  assign n5919 = ~n5911 & n5918;
  assign n5920 = n5911 & ~n5918;
  assign n5921 = ~n5919 & ~n5920;
  assign n5922 = A904  & A905 ;
  assign n5923 = A906  & ~n5916;
  assign n5924 = ~n5922 & ~n5923;
  assign n5925 = A901  & A902 ;
  assign n5926 = A903  & ~n5909;
  assign n5927 = ~n5925 & ~n5926;
  assign n5928 = ~n5924 & n5927;
  assign n5929 = n5924 & ~n5927;
  assign n5930 = ~n5928 & ~n5929;
  assign n5931 = ~n5911 & ~n5918;
  assign n5932 = ~n5930 & n5931;
  assign n5933 = ~n5924 & ~n5927;
  assign n5934 = ~n5932 & ~n5933;
  assign n5935 = ~n5928 & n5931;
  assign n5936 = ~n5929 & n5935;
  assign n5937 = ~n5930 & ~n5931;
  assign n5938 = ~n5936 & ~n5937;
  assign n5939 = ~n5934 & ~n5938;
  assign n5940 = ~n5921 & ~n5939;
  assign n5941 = ~A895  & A896 ;
  assign n5942 = A895  & ~A896 ;
  assign n5943 = A897  & ~n5942;
  assign n5944 = ~n5941 & n5943;
  assign n5945 = ~n5941 & ~n5942;
  assign n5946 = ~A897  & ~n5945;
  assign n5947 = ~n5944 & ~n5946;
  assign n5948 = ~A898  & A899 ;
  assign n5949 = A898  & ~A899 ;
  assign n5950 = A900  & ~n5949;
  assign n5951 = ~n5948 & n5950;
  assign n5952 = ~n5948 & ~n5949;
  assign n5953 = ~A900  & ~n5952;
  assign n5954 = ~n5951 & ~n5953;
  assign n5955 = ~n5947 & n5954;
  assign n5956 = n5947 & ~n5954;
  assign n5957 = ~n5955 & ~n5956;
  assign n5958 = A898  & A899 ;
  assign n5959 = A900  & ~n5952;
  assign n5960 = ~n5958 & ~n5959;
  assign n5961 = A895  & A896 ;
  assign n5962 = A897  & ~n5945;
  assign n5963 = ~n5961 & ~n5962;
  assign n5964 = ~n5960 & n5963;
  assign n5965 = n5960 & ~n5963;
  assign n5966 = ~n5964 & ~n5965;
  assign n5967 = ~n5947 & ~n5954;
  assign n5968 = ~n5966 & n5967;
  assign n5969 = ~n5960 & ~n5963;
  assign n5970 = ~n5968 & ~n5969;
  assign n5971 = ~n5964 & n5967;
  assign n5972 = ~n5965 & n5971;
  assign n5973 = ~n5966 & ~n5967;
  assign n5974 = ~n5972 & ~n5973;
  assign n5975 = ~n5970 & ~n5974;
  assign n5976 = ~n5957 & ~n5975;
  assign n5977 = ~n5940 & n5976;
  assign n5978 = n5940 & ~n5976;
  assign n5979 = ~n5977 & ~n5978;
  assign n5980 = ~n5904 & n5979;
  assign n5981 = n5904 & ~n5979;
  assign n5982 = ~n5980 & ~n5981;
  assign n5983 = ~n5829 & n5982;
  assign n5984 = n5829 & ~n5982;
  assign n5985 = ~n5983 & ~n5984;
  assign n5986 = ~A889  & A890 ;
  assign n5987 = A889  & ~A890 ;
  assign n5988 = A891  & ~n5987;
  assign n5989 = ~n5986 & n5988;
  assign n5990 = ~n5986 & ~n5987;
  assign n5991 = ~A891  & ~n5990;
  assign n5992 = ~n5989 & ~n5991;
  assign n5993 = ~A892  & A893 ;
  assign n5994 = A892  & ~A893 ;
  assign n5995 = A894  & ~n5994;
  assign n5996 = ~n5993 & n5995;
  assign n5997 = ~n5993 & ~n5994;
  assign n5998 = ~A894  & ~n5997;
  assign n5999 = ~n5996 & ~n5998;
  assign n6000 = ~n5992 & n5999;
  assign n6001 = n5992 & ~n5999;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = A892  & A893 ;
  assign n6004 = A894  & ~n5997;
  assign n6005 = ~n6003 & ~n6004;
  assign n6006 = A889  & A890 ;
  assign n6007 = A891  & ~n5990;
  assign n6008 = ~n6006 & ~n6007;
  assign n6009 = ~n6005 & n6008;
  assign n6010 = n6005 & ~n6008;
  assign n6011 = ~n6009 & ~n6010;
  assign n6012 = ~n5992 & ~n5999;
  assign n6013 = ~n6011 & n6012;
  assign n6014 = ~n6005 & ~n6008;
  assign n6015 = ~n6013 & ~n6014;
  assign n6016 = ~n6009 & n6012;
  assign n6017 = ~n6010 & n6016;
  assign n6018 = ~n6011 & ~n6012;
  assign n6019 = ~n6017 & ~n6018;
  assign n6020 = ~n6015 & ~n6019;
  assign n6021 = ~n6002 & ~n6020;
  assign n6022 = ~A883  & A884 ;
  assign n6023 = A883  & ~A884 ;
  assign n6024 = A885  & ~n6023;
  assign n6025 = ~n6022 & n6024;
  assign n6026 = ~n6022 & ~n6023;
  assign n6027 = ~A885  & ~n6026;
  assign n6028 = ~n6025 & ~n6027;
  assign n6029 = ~A886  & A887 ;
  assign n6030 = A886  & ~A887 ;
  assign n6031 = A888  & ~n6030;
  assign n6032 = ~n6029 & n6031;
  assign n6033 = ~n6029 & ~n6030;
  assign n6034 = ~A888  & ~n6033;
  assign n6035 = ~n6032 & ~n6034;
  assign n6036 = ~n6028 & n6035;
  assign n6037 = n6028 & ~n6035;
  assign n6038 = ~n6036 & ~n6037;
  assign n6039 = A886  & A887 ;
  assign n6040 = A888  & ~n6033;
  assign n6041 = ~n6039 & ~n6040;
  assign n6042 = A883  & A884 ;
  assign n6043 = A885  & ~n6026;
  assign n6044 = ~n6042 & ~n6043;
  assign n6045 = ~n6041 & n6044;
  assign n6046 = n6041 & ~n6044;
  assign n6047 = ~n6045 & ~n6046;
  assign n6048 = ~n6028 & ~n6035;
  assign n6049 = ~n6047 & n6048;
  assign n6050 = ~n6041 & ~n6044;
  assign n6051 = ~n6049 & ~n6050;
  assign n6052 = ~n6045 & n6048;
  assign n6053 = ~n6046 & n6052;
  assign n6054 = ~n6047 & ~n6048;
  assign n6055 = ~n6053 & ~n6054;
  assign n6056 = ~n6051 & ~n6055;
  assign n6057 = ~n6038 & ~n6056;
  assign n6058 = ~n6021 & n6057;
  assign n6059 = n6021 & ~n6057;
  assign n6060 = ~n6058 & ~n6059;
  assign n6061 = ~A877  & A878 ;
  assign n6062 = A877  & ~A878 ;
  assign n6063 = A879  & ~n6062;
  assign n6064 = ~n6061 & n6063;
  assign n6065 = ~n6061 & ~n6062;
  assign n6066 = ~A879  & ~n6065;
  assign n6067 = ~n6064 & ~n6066;
  assign n6068 = ~A880  & A881 ;
  assign n6069 = A880  & ~A881 ;
  assign n6070 = A882  & ~n6069;
  assign n6071 = ~n6068 & n6070;
  assign n6072 = ~n6068 & ~n6069;
  assign n6073 = ~A882  & ~n6072;
  assign n6074 = ~n6071 & ~n6073;
  assign n6075 = ~n6067 & n6074;
  assign n6076 = n6067 & ~n6074;
  assign n6077 = ~n6075 & ~n6076;
  assign n6078 = A880  & A881 ;
  assign n6079 = A882  & ~n6072;
  assign n6080 = ~n6078 & ~n6079;
  assign n6081 = A877  & A878 ;
  assign n6082 = A879  & ~n6065;
  assign n6083 = ~n6081 & ~n6082;
  assign n6084 = ~n6080 & n6083;
  assign n6085 = n6080 & ~n6083;
  assign n6086 = ~n6084 & ~n6085;
  assign n6087 = ~n6067 & ~n6074;
  assign n6088 = ~n6086 & n6087;
  assign n6089 = ~n6080 & ~n6083;
  assign n6090 = ~n6088 & ~n6089;
  assign n6091 = ~n6084 & n6087;
  assign n6092 = ~n6085 & n6091;
  assign n6093 = ~n6086 & ~n6087;
  assign n6094 = ~n6092 & ~n6093;
  assign n6095 = ~n6090 & ~n6094;
  assign n6096 = ~n6077 & ~n6095;
  assign n6097 = ~A871  & A872 ;
  assign n6098 = A871  & ~A872 ;
  assign n6099 = A873  & ~n6098;
  assign n6100 = ~n6097 & n6099;
  assign n6101 = ~n6097 & ~n6098;
  assign n6102 = ~A873  & ~n6101;
  assign n6103 = ~n6100 & ~n6102;
  assign n6104 = ~A874  & A875 ;
  assign n6105 = A874  & ~A875 ;
  assign n6106 = A876  & ~n6105;
  assign n6107 = ~n6104 & n6106;
  assign n6108 = ~n6104 & ~n6105;
  assign n6109 = ~A876  & ~n6108;
  assign n6110 = ~n6107 & ~n6109;
  assign n6111 = ~n6103 & n6110;
  assign n6112 = n6103 & ~n6110;
  assign n6113 = ~n6111 & ~n6112;
  assign n6114 = A874  & A875 ;
  assign n6115 = A876  & ~n6108;
  assign n6116 = ~n6114 & ~n6115;
  assign n6117 = A871  & A872 ;
  assign n6118 = A873  & ~n6101;
  assign n6119 = ~n6117 & ~n6118;
  assign n6120 = ~n6116 & n6119;
  assign n6121 = n6116 & ~n6119;
  assign n6122 = ~n6120 & ~n6121;
  assign n6123 = ~n6103 & ~n6110;
  assign n6124 = ~n6122 & n6123;
  assign n6125 = ~n6116 & ~n6119;
  assign n6126 = ~n6124 & ~n6125;
  assign n6127 = ~n6120 & n6123;
  assign n6128 = ~n6121 & n6127;
  assign n6129 = ~n6122 & ~n6123;
  assign n6130 = ~n6128 & ~n6129;
  assign n6131 = ~n6126 & ~n6130;
  assign n6132 = ~n6113 & ~n6131;
  assign n6133 = ~n6096 & n6132;
  assign n6134 = n6096 & ~n6132;
  assign n6135 = ~n6133 & ~n6134;
  assign n6136 = ~n6060 & n6135;
  assign n6137 = n6060 & ~n6135;
  assign n6138 = ~n6136 & ~n6137;
  assign n6139 = ~A865  & A866 ;
  assign n6140 = A865  & ~A866 ;
  assign n6141 = A867  & ~n6140;
  assign n6142 = ~n6139 & n6141;
  assign n6143 = ~n6139 & ~n6140;
  assign n6144 = ~A867  & ~n6143;
  assign n6145 = ~n6142 & ~n6144;
  assign n6146 = ~A868  & A869 ;
  assign n6147 = A868  & ~A869 ;
  assign n6148 = A870  & ~n6147;
  assign n6149 = ~n6146 & n6148;
  assign n6150 = ~n6146 & ~n6147;
  assign n6151 = ~A870  & ~n6150;
  assign n6152 = ~n6149 & ~n6151;
  assign n6153 = ~n6145 & n6152;
  assign n6154 = n6145 & ~n6152;
  assign n6155 = ~n6153 & ~n6154;
  assign n6156 = A868  & A869 ;
  assign n6157 = A870  & ~n6150;
  assign n6158 = ~n6156 & ~n6157;
  assign n6159 = A865  & A866 ;
  assign n6160 = A867  & ~n6143;
  assign n6161 = ~n6159 & ~n6160;
  assign n6162 = ~n6158 & n6161;
  assign n6163 = n6158 & ~n6161;
  assign n6164 = ~n6162 & ~n6163;
  assign n6165 = ~n6145 & ~n6152;
  assign n6166 = ~n6164 & n6165;
  assign n6167 = ~n6158 & ~n6161;
  assign n6168 = ~n6166 & ~n6167;
  assign n6169 = ~n6162 & n6165;
  assign n6170 = ~n6163 & n6169;
  assign n6171 = ~n6164 & ~n6165;
  assign n6172 = ~n6170 & ~n6171;
  assign n6173 = ~n6168 & ~n6172;
  assign n6174 = ~n6155 & ~n6173;
  assign n6175 = ~A859  & A860 ;
  assign n6176 = A859  & ~A860 ;
  assign n6177 = A861  & ~n6176;
  assign n6178 = ~n6175 & n6177;
  assign n6179 = ~n6175 & ~n6176;
  assign n6180 = ~A861  & ~n6179;
  assign n6181 = ~n6178 & ~n6180;
  assign n6182 = ~A862  & A863 ;
  assign n6183 = A862  & ~A863 ;
  assign n6184 = A864  & ~n6183;
  assign n6185 = ~n6182 & n6184;
  assign n6186 = ~n6182 & ~n6183;
  assign n6187 = ~A864  & ~n6186;
  assign n6188 = ~n6185 & ~n6187;
  assign n6189 = ~n6181 & n6188;
  assign n6190 = n6181 & ~n6188;
  assign n6191 = ~n6189 & ~n6190;
  assign n6192 = A862  & A863 ;
  assign n6193 = A864  & ~n6186;
  assign n6194 = ~n6192 & ~n6193;
  assign n6195 = A859  & A860 ;
  assign n6196 = A861  & ~n6179;
  assign n6197 = ~n6195 & ~n6196;
  assign n6198 = ~n6194 & n6197;
  assign n6199 = n6194 & ~n6197;
  assign n6200 = ~n6198 & ~n6199;
  assign n6201 = ~n6181 & ~n6188;
  assign n6202 = ~n6200 & n6201;
  assign n6203 = ~n6194 & ~n6197;
  assign n6204 = ~n6202 & ~n6203;
  assign n6205 = ~n6198 & n6201;
  assign n6206 = ~n6199 & n6205;
  assign n6207 = ~n6200 & ~n6201;
  assign n6208 = ~n6206 & ~n6207;
  assign n6209 = ~n6204 & ~n6208;
  assign n6210 = ~n6191 & ~n6209;
  assign n6211 = ~n6174 & n6210;
  assign n6212 = n6174 & ~n6210;
  assign n6213 = ~n6211 & ~n6212;
  assign n6214 = ~A853  & A854 ;
  assign n6215 = A853  & ~A854 ;
  assign n6216 = A855  & ~n6215;
  assign n6217 = ~n6214 & n6216;
  assign n6218 = ~n6214 & ~n6215;
  assign n6219 = ~A855  & ~n6218;
  assign n6220 = ~n6217 & ~n6219;
  assign n6221 = ~A856  & A857 ;
  assign n6222 = A856  & ~A857 ;
  assign n6223 = A858  & ~n6222;
  assign n6224 = ~n6221 & n6223;
  assign n6225 = ~n6221 & ~n6222;
  assign n6226 = ~A858  & ~n6225;
  assign n6227 = ~n6224 & ~n6226;
  assign n6228 = ~n6220 & n6227;
  assign n6229 = n6220 & ~n6227;
  assign n6230 = ~n6228 & ~n6229;
  assign n6231 = A856  & A857 ;
  assign n6232 = A858  & ~n6225;
  assign n6233 = ~n6231 & ~n6232;
  assign n6234 = A853  & A854 ;
  assign n6235 = A855  & ~n6218;
  assign n6236 = ~n6234 & ~n6235;
  assign n6237 = ~n6233 & n6236;
  assign n6238 = n6233 & ~n6236;
  assign n6239 = ~n6237 & ~n6238;
  assign n6240 = ~n6220 & ~n6227;
  assign n6241 = ~n6239 & n6240;
  assign n6242 = ~n6233 & ~n6236;
  assign n6243 = ~n6241 & ~n6242;
  assign n6244 = ~n6237 & n6240;
  assign n6245 = ~n6238 & n6244;
  assign n6246 = ~n6239 & ~n6240;
  assign n6247 = ~n6245 & ~n6246;
  assign n6248 = ~n6243 & ~n6247;
  assign n6249 = ~n6230 & ~n6248;
  assign n6250 = ~A847  & A848 ;
  assign n6251 = A847  & ~A848 ;
  assign n6252 = A849  & ~n6251;
  assign n6253 = ~n6250 & n6252;
  assign n6254 = ~n6250 & ~n6251;
  assign n6255 = ~A849  & ~n6254;
  assign n6256 = ~n6253 & ~n6255;
  assign n6257 = ~A850  & A851 ;
  assign n6258 = A850  & ~A851 ;
  assign n6259 = A852  & ~n6258;
  assign n6260 = ~n6257 & n6259;
  assign n6261 = ~n6257 & ~n6258;
  assign n6262 = ~A852  & ~n6261;
  assign n6263 = ~n6260 & ~n6262;
  assign n6264 = ~n6256 & n6263;
  assign n6265 = n6256 & ~n6263;
  assign n6266 = ~n6264 & ~n6265;
  assign n6267 = A850  & A851 ;
  assign n6268 = A852  & ~n6261;
  assign n6269 = ~n6267 & ~n6268;
  assign n6270 = A847  & A848 ;
  assign n6271 = A849  & ~n6254;
  assign n6272 = ~n6270 & ~n6271;
  assign n6273 = ~n6269 & n6272;
  assign n6274 = n6269 & ~n6272;
  assign n6275 = ~n6273 & ~n6274;
  assign n6276 = ~n6256 & ~n6263;
  assign n6277 = ~n6275 & n6276;
  assign n6278 = ~n6269 & ~n6272;
  assign n6279 = ~n6277 & ~n6278;
  assign n6280 = ~n6273 & n6276;
  assign n6281 = ~n6274 & n6280;
  assign n6282 = ~n6275 & ~n6276;
  assign n6283 = ~n6281 & ~n6282;
  assign n6284 = ~n6279 & ~n6283;
  assign n6285 = ~n6266 & ~n6284;
  assign n6286 = ~n6249 & n6285;
  assign n6287 = n6249 & ~n6285;
  assign n6288 = ~n6286 & ~n6287;
  assign n6289 = ~n6213 & n6288;
  assign n6290 = n6213 & ~n6288;
  assign n6291 = ~n6289 & ~n6290;
  assign n6292 = ~n6138 & n6291;
  assign n6293 = n6138 & ~n6291;
  assign n6294 = ~n6292 & ~n6293;
  assign n6295 = ~n5985 & n6294;
  assign n6296 = n5985 & ~n6294;
  assign n6297 = ~n6295 & ~n6296;
  assign n6298 = ~n5676 & ~n6297;
  assign n6299 = ~n5672 & n6298;
  assign n6300 = ~n5667 & n6299;
  assign n6301 = ~n5667 & ~n5672;
  assign n6302 = ~n6298 & ~n6301;
  assign n6303 = ~n6300 & ~n6302;
  assign n6304 = ~n5882 & ~n5895;
  assign n6305 = ~n5899 & ~n6304;
  assign n6306 = ~n5846 & ~n5882;
  assign n6307 = ~n5864 & n6306;
  assign n6308 = ~n5900 & n6307;
  assign n6309 = ~n5846 & ~n5859;
  assign n6310 = ~n5863 & ~n6309;
  assign n6311 = ~n6308 & ~n6310;
  assign n6312 = ~n5863 & n6306;
  assign n6313 = ~n5864 & n6312;
  assign n6314 = ~n5900 & ~n6309;
  assign n6315 = n6313 & n6314;
  assign n6316 = ~n6311 & ~n6315;
  assign n6317 = n6305 & ~n6316;
  assign n6318 = ~n6308 & n6310;
  assign n6319 = n6308 & ~n6310;
  assign n6320 = ~n6318 & ~n6319;
  assign n6321 = ~n6305 & ~n6320;
  assign n6322 = ~n5904 & ~n5979;
  assign n6323 = ~n6321 & n6322;
  assign n6324 = ~n6317 & n6323;
  assign n6325 = ~n6317 & ~n6321;
  assign n6326 = ~n6322 & ~n6325;
  assign n6327 = ~n6324 & ~n6326;
  assign n6328 = ~n5957 & ~n5970;
  assign n6329 = ~n5974 & ~n6328;
  assign n6330 = ~n5921 & ~n5957;
  assign n6331 = ~n5939 & n6330;
  assign n6332 = ~n5975 & n6331;
  assign n6333 = ~n5921 & ~n5934;
  assign n6334 = ~n5938 & ~n6333;
  assign n6335 = ~n6332 & n6334;
  assign n6336 = n6332 & ~n6334;
  assign n6337 = ~n6335 & ~n6336;
  assign n6338 = ~n6329 & ~n6337;
  assign n6339 = ~n6332 & ~n6334;
  assign n6340 = ~n5938 & n6330;
  assign n6341 = ~n5939 & n6340;
  assign n6342 = ~n5975 & ~n6333;
  assign n6343 = n6341 & n6342;
  assign n6344 = ~n6339 & ~n6343;
  assign n6345 = n6329 & ~n6344;
  assign n6346 = ~n6338 & ~n6345;
  assign n6347 = ~n6327 & n6346;
  assign n6348 = ~n6321 & ~n6322;
  assign n6349 = ~n6317 & n6348;
  assign n6350 = n6322 & ~n6325;
  assign n6351 = ~n6349 & ~n6350;
  assign n6352 = ~n6346 & ~n6351;
  assign n6353 = ~n6347 & ~n6352;
  assign n6354 = ~n5804 & ~n5817;
  assign n6355 = ~n5821 & ~n6354;
  assign n6356 = ~n5768 & ~n5804;
  assign n6357 = ~n5786 & n6356;
  assign n6358 = ~n5822 & n6357;
  assign n6359 = ~n5768 & ~n5781;
  assign n6360 = ~n5785 & ~n6359;
  assign n6361 = ~n6358 & n6360;
  assign n6362 = n6358 & ~n6360;
  assign n6363 = ~n6361 & ~n6362;
  assign n6364 = ~n6355 & ~n6363;
  assign n6365 = ~n6358 & ~n6360;
  assign n6366 = ~n5785 & n6356;
  assign n6367 = ~n5786 & n6366;
  assign n6368 = ~n5822 & ~n6359;
  assign n6369 = n6367 & n6368;
  assign n6370 = ~n6365 & ~n6369;
  assign n6371 = n6355 & ~n6370;
  assign n6372 = ~n6364 & ~n6371;
  assign n6373 = ~n5729 & ~n5742;
  assign n6374 = ~n5746 & ~n6373;
  assign n6375 = ~n5693 & ~n5729;
  assign n6376 = ~n5711 & n6375;
  assign n6377 = ~n5747 & n6376;
  assign n6378 = ~n5693 & ~n5706;
  assign n6379 = ~n5710 & ~n6378;
  assign n6380 = ~n6377 & ~n6379;
  assign n6381 = ~n5710 & n6375;
  assign n6382 = ~n5711 & n6381;
  assign n6383 = ~n5747 & ~n6378;
  assign n6384 = n6382 & n6383;
  assign n6385 = ~n6380 & ~n6384;
  assign n6386 = n6374 & ~n6385;
  assign n6387 = ~n6377 & n6379;
  assign n6388 = n6377 & ~n6379;
  assign n6389 = ~n6387 & ~n6388;
  assign n6390 = ~n6374 & ~n6389;
  assign n6391 = ~n5751 & ~n5826;
  assign n6392 = ~n6390 & ~n6391;
  assign n6393 = ~n6386 & n6392;
  assign n6394 = ~n6386 & ~n6390;
  assign n6395 = n6391 & ~n6394;
  assign n6396 = ~n6393 & ~n6395;
  assign n6397 = ~n6372 & ~n6396;
  assign n6398 = ~n6390 & n6391;
  assign n6399 = ~n6386 & n6398;
  assign n6400 = ~n6391 & ~n6394;
  assign n6401 = ~n6399 & ~n6400;
  assign n6402 = n6372 & ~n6401;
  assign n6403 = ~n5829 & ~n5982;
  assign n6404 = ~n6402 & ~n6403;
  assign n6405 = ~n6397 & n6404;
  assign n6406 = ~n6397 & ~n6402;
  assign n6407 = n6403 & ~n6406;
  assign n6408 = ~n6405 & ~n6407;
  assign n6409 = ~n6353 & ~n6408;
  assign n6410 = ~n6402 & n6403;
  assign n6411 = ~n6397 & n6410;
  assign n6412 = ~n6403 & ~n6406;
  assign n6413 = ~n6411 & ~n6412;
  assign n6414 = n6353 & ~n6413;
  assign n6415 = ~n5985 & ~n6294;
  assign n6416 = ~n6414 & n6415;
  assign n6417 = ~n6409 & n6416;
  assign n6418 = ~n6409 & ~n6414;
  assign n6419 = ~n6415 & ~n6418;
  assign n6420 = ~n6417 & ~n6419;
  assign n6421 = ~n6113 & ~n6126;
  assign n6422 = ~n6130 & ~n6421;
  assign n6423 = ~n6077 & ~n6113;
  assign n6424 = ~n6095 & n6423;
  assign n6425 = ~n6131 & n6424;
  assign n6426 = ~n6077 & ~n6090;
  assign n6427 = ~n6094 & ~n6426;
  assign n6428 = ~n6425 & n6427;
  assign n6429 = n6425 & ~n6427;
  assign n6430 = ~n6428 & ~n6429;
  assign n6431 = ~n6422 & ~n6430;
  assign n6432 = ~n6425 & ~n6427;
  assign n6433 = ~n6094 & n6423;
  assign n6434 = ~n6095 & n6433;
  assign n6435 = ~n6131 & ~n6426;
  assign n6436 = n6434 & n6435;
  assign n6437 = ~n6432 & ~n6436;
  assign n6438 = n6422 & ~n6437;
  assign n6439 = ~n6431 & ~n6438;
  assign n6440 = ~n6038 & ~n6051;
  assign n6441 = ~n6055 & ~n6440;
  assign n6442 = ~n6002 & ~n6038;
  assign n6443 = ~n6020 & n6442;
  assign n6444 = ~n6056 & n6443;
  assign n6445 = ~n6002 & ~n6015;
  assign n6446 = ~n6019 & ~n6445;
  assign n6447 = ~n6444 & ~n6446;
  assign n6448 = ~n6019 & n6442;
  assign n6449 = ~n6020 & n6448;
  assign n6450 = ~n6056 & ~n6445;
  assign n6451 = n6449 & n6450;
  assign n6452 = ~n6447 & ~n6451;
  assign n6453 = n6441 & ~n6452;
  assign n6454 = ~n6444 & n6446;
  assign n6455 = n6444 & ~n6446;
  assign n6456 = ~n6454 & ~n6455;
  assign n6457 = ~n6441 & ~n6456;
  assign n6458 = ~n6060 & ~n6135;
  assign n6459 = ~n6457 & ~n6458;
  assign n6460 = ~n6453 & n6459;
  assign n6461 = ~n6453 & ~n6457;
  assign n6462 = n6458 & ~n6461;
  assign n6463 = ~n6460 & ~n6462;
  assign n6464 = ~n6439 & ~n6463;
  assign n6465 = ~n6457 & n6458;
  assign n6466 = ~n6453 & n6465;
  assign n6467 = ~n6458 & ~n6461;
  assign n6468 = ~n6466 & ~n6467;
  assign n6469 = n6439 & ~n6468;
  assign n6470 = ~n6138 & ~n6291;
  assign n6471 = ~n6469 & n6470;
  assign n6472 = ~n6464 & n6471;
  assign n6473 = ~n6464 & ~n6469;
  assign n6474 = ~n6470 & ~n6473;
  assign n6475 = ~n6472 & ~n6474;
  assign n6476 = ~n6191 & ~n6204;
  assign n6477 = ~n6208 & ~n6476;
  assign n6478 = ~n6155 & ~n6191;
  assign n6479 = ~n6173 & n6478;
  assign n6480 = ~n6209 & n6479;
  assign n6481 = ~n6155 & ~n6168;
  assign n6482 = ~n6172 & ~n6481;
  assign n6483 = ~n6480 & ~n6482;
  assign n6484 = ~n6172 & n6478;
  assign n6485 = ~n6173 & n6484;
  assign n6486 = ~n6209 & ~n6481;
  assign n6487 = n6485 & n6486;
  assign n6488 = ~n6483 & ~n6487;
  assign n6489 = n6477 & ~n6488;
  assign n6490 = ~n6480 & n6482;
  assign n6491 = n6480 & ~n6482;
  assign n6492 = ~n6490 & ~n6491;
  assign n6493 = ~n6477 & ~n6492;
  assign n6494 = ~n6213 & ~n6288;
  assign n6495 = ~n6493 & n6494;
  assign n6496 = ~n6489 & n6495;
  assign n6497 = ~n6489 & ~n6493;
  assign n6498 = ~n6494 & ~n6497;
  assign n6499 = ~n6496 & ~n6498;
  assign n6500 = ~n6266 & ~n6279;
  assign n6501 = ~n6283 & ~n6500;
  assign n6502 = ~n6230 & ~n6266;
  assign n6503 = ~n6248 & n6502;
  assign n6504 = ~n6284 & n6503;
  assign n6505 = ~n6230 & ~n6243;
  assign n6506 = ~n6247 & ~n6505;
  assign n6507 = ~n6504 & n6506;
  assign n6508 = n6504 & ~n6506;
  assign n6509 = ~n6507 & ~n6508;
  assign n6510 = ~n6501 & ~n6509;
  assign n6511 = ~n6504 & ~n6506;
  assign n6512 = ~n6247 & n6502;
  assign n6513 = ~n6248 & n6512;
  assign n6514 = ~n6284 & ~n6505;
  assign n6515 = n6513 & n6514;
  assign n6516 = ~n6511 & ~n6515;
  assign n6517 = n6501 & ~n6516;
  assign n6518 = ~n6510 & ~n6517;
  assign n6519 = ~n6499 & n6518;
  assign n6520 = ~n6493 & ~n6494;
  assign n6521 = ~n6489 & n6520;
  assign n6522 = n6494 & ~n6497;
  assign n6523 = ~n6521 & ~n6522;
  assign n6524 = ~n6518 & ~n6523;
  assign n6525 = ~n6519 & ~n6524;
  assign n6526 = ~n6475 & n6525;
  assign n6527 = ~n6469 & ~n6470;
  assign n6528 = ~n6464 & n6527;
  assign n6529 = n6470 & ~n6473;
  assign n6530 = ~n6528 & ~n6529;
  assign n6531 = ~n6525 & ~n6530;
  assign n6532 = ~n6526 & ~n6531;
  assign n6533 = ~n6420 & n6532;
  assign n6534 = ~n6414 & ~n6415;
  assign n6535 = ~n6409 & n6534;
  assign n6536 = n6415 & ~n6418;
  assign n6537 = ~n6535 & ~n6536;
  assign n6538 = ~n6532 & ~n6537;
  assign n6539 = ~n6533 & ~n6538;
  assign n6540 = ~n6303 & n6539;
  assign n6541 = ~n5672 & ~n6298;
  assign n6542 = ~n5667 & n6541;
  assign n6543 = n6298 & ~n6301;
  assign n6544 = ~n6542 & ~n6543;
  assign n6545 = ~n6539 & ~n6544;
  assign n6546 = ~n6540 & ~n6545;
  assign n6547 = A202  & A203 ;
  assign n6548 = A202  & ~A203 ;
  assign n6549 = ~A202  & A203 ;
  assign n6550 = ~n6548 & ~n6549;
  assign n6551 = A204  & ~n6550;
  assign n6552 = ~n6547 & ~n6551;
  assign n6553 = A199  & A200 ;
  assign n6554 = A199  & ~A200 ;
  assign n6555 = ~A199  & A200 ;
  assign n6556 = ~n6554 & ~n6555;
  assign n6557 = A201  & ~n6556;
  assign n6558 = ~n6553 & ~n6557;
  assign n6559 = n6552 & ~n6558;
  assign n6560 = ~n6552 & n6558;
  assign n6561 = A201  & ~n6554;
  assign n6562 = ~n6555 & n6561;
  assign n6563 = ~A201  & ~n6556;
  assign n6564 = ~n6562 & ~n6563;
  assign n6565 = A204  & ~n6548;
  assign n6566 = ~n6549 & n6565;
  assign n6567 = ~A204  & ~n6550;
  assign n6568 = ~n6566 & ~n6567;
  assign n6569 = ~n6564 & ~n6568;
  assign n6570 = ~n6560 & n6569;
  assign n6571 = ~n6559 & n6570;
  assign n6572 = ~n6559 & ~n6560;
  assign n6573 = ~n6569 & ~n6572;
  assign n6574 = ~n6571 & ~n6573;
  assign n6575 = ~n6564 & n6568;
  assign n6576 = n6564 & ~n6568;
  assign n6577 = ~n6575 & ~n6576;
  assign n6578 = n6569 & ~n6572;
  assign n6579 = ~n6552 & ~n6558;
  assign n6580 = ~n6578 & ~n6579;
  assign n6581 = ~n6577 & ~n6580;
  assign n6582 = ~n6574 & ~n6581;
  assign n6583 = ~n6574 & ~n6580;
  assign n6584 = A208  & A209 ;
  assign n6585 = A208  & ~A209 ;
  assign n6586 = ~A208  & A209 ;
  assign n6587 = ~n6585 & ~n6586;
  assign n6588 = A210  & ~n6587;
  assign n6589 = ~n6584 & ~n6588;
  assign n6590 = A205  & A206 ;
  assign n6591 = A205  & ~A206 ;
  assign n6592 = ~A205  & A206 ;
  assign n6593 = ~n6591 & ~n6592;
  assign n6594 = A207  & ~n6593;
  assign n6595 = ~n6590 & ~n6594;
  assign n6596 = ~n6589 & n6595;
  assign n6597 = n6589 & ~n6595;
  assign n6598 = ~n6596 & ~n6597;
  assign n6599 = A207  & ~n6591;
  assign n6600 = ~n6592 & n6599;
  assign n6601 = ~A207  & ~n6593;
  assign n6602 = ~n6600 & ~n6601;
  assign n6603 = A210  & ~n6585;
  assign n6604 = ~n6586 & n6603;
  assign n6605 = ~A210  & ~n6587;
  assign n6606 = ~n6604 & ~n6605;
  assign n6607 = ~n6602 & ~n6606;
  assign n6608 = ~n6598 & n6607;
  assign n6609 = ~n6589 & ~n6595;
  assign n6610 = ~n6608 & ~n6609;
  assign n6611 = ~n6596 & n6607;
  assign n6612 = ~n6597 & n6611;
  assign n6613 = ~n6598 & ~n6607;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = ~n6610 & ~n6614;
  assign n6616 = ~n6602 & n6606;
  assign n6617 = n6602 & ~n6606;
  assign n6618 = ~n6616 & ~n6617;
  assign n6619 = ~n6577 & ~n6618;
  assign n6620 = ~n6615 & n6619;
  assign n6621 = ~n6583 & n6620;
  assign n6622 = ~n6610 & ~n6618;
  assign n6623 = ~n6614 & ~n6622;
  assign n6624 = ~n6621 & n6623;
  assign n6625 = n6621 & ~n6623;
  assign n6626 = ~n6624 & ~n6625;
  assign n6627 = ~n6582 & ~n6626;
  assign n6628 = ~n6621 & ~n6623;
  assign n6629 = ~n6614 & n6619;
  assign n6630 = ~n6615 & n6629;
  assign n6631 = ~n6583 & ~n6622;
  assign n6632 = n6630 & n6631;
  assign n6633 = ~n6628 & ~n6632;
  assign n6634 = n6582 & ~n6633;
  assign n6635 = ~n6627 & ~n6634;
  assign n6636 = A214  & A215 ;
  assign n6637 = A214  & ~A215 ;
  assign n6638 = ~A214  & A215 ;
  assign n6639 = ~n6637 & ~n6638;
  assign n6640 = A216  & ~n6639;
  assign n6641 = ~n6636 & ~n6640;
  assign n6642 = A211  & A212 ;
  assign n6643 = A211  & ~A212 ;
  assign n6644 = ~A211  & A212 ;
  assign n6645 = ~n6643 & ~n6644;
  assign n6646 = A213  & ~n6645;
  assign n6647 = ~n6642 & ~n6646;
  assign n6648 = n6641 & ~n6647;
  assign n6649 = ~n6641 & n6647;
  assign n6650 = A213  & ~n6643;
  assign n6651 = ~n6644 & n6650;
  assign n6652 = ~A213  & ~n6645;
  assign n6653 = ~n6651 & ~n6652;
  assign n6654 = A216  & ~n6637;
  assign n6655 = ~n6638 & n6654;
  assign n6656 = ~A216  & ~n6639;
  assign n6657 = ~n6655 & ~n6656;
  assign n6658 = ~n6653 & ~n6657;
  assign n6659 = ~n6649 & n6658;
  assign n6660 = ~n6648 & n6659;
  assign n6661 = ~n6648 & ~n6649;
  assign n6662 = ~n6658 & ~n6661;
  assign n6663 = ~n6660 & ~n6662;
  assign n6664 = ~n6653 & n6657;
  assign n6665 = n6653 & ~n6657;
  assign n6666 = ~n6664 & ~n6665;
  assign n6667 = n6658 & ~n6661;
  assign n6668 = ~n6641 & ~n6647;
  assign n6669 = ~n6667 & ~n6668;
  assign n6670 = ~n6666 & ~n6669;
  assign n6671 = ~n6663 & ~n6670;
  assign n6672 = ~n6663 & ~n6669;
  assign n6673 = A220  & A221 ;
  assign n6674 = A220  & ~A221 ;
  assign n6675 = ~A220  & A221 ;
  assign n6676 = ~n6674 & ~n6675;
  assign n6677 = A222  & ~n6676;
  assign n6678 = ~n6673 & ~n6677;
  assign n6679 = A217  & A218 ;
  assign n6680 = A217  & ~A218 ;
  assign n6681 = ~A217  & A218 ;
  assign n6682 = ~n6680 & ~n6681;
  assign n6683 = A219  & ~n6682;
  assign n6684 = ~n6679 & ~n6683;
  assign n6685 = ~n6678 & n6684;
  assign n6686 = n6678 & ~n6684;
  assign n6687 = ~n6685 & ~n6686;
  assign n6688 = A219  & ~n6680;
  assign n6689 = ~n6681 & n6688;
  assign n6690 = ~A219  & ~n6682;
  assign n6691 = ~n6689 & ~n6690;
  assign n6692 = A222  & ~n6674;
  assign n6693 = ~n6675 & n6692;
  assign n6694 = ~A222  & ~n6676;
  assign n6695 = ~n6693 & ~n6694;
  assign n6696 = ~n6691 & ~n6695;
  assign n6697 = ~n6687 & n6696;
  assign n6698 = ~n6678 & ~n6684;
  assign n6699 = ~n6697 & ~n6698;
  assign n6700 = ~n6685 & n6696;
  assign n6701 = ~n6686 & n6700;
  assign n6702 = ~n6687 & ~n6696;
  assign n6703 = ~n6701 & ~n6702;
  assign n6704 = ~n6699 & ~n6703;
  assign n6705 = ~n6691 & n6695;
  assign n6706 = n6691 & ~n6695;
  assign n6707 = ~n6705 & ~n6706;
  assign n6708 = ~n6666 & ~n6707;
  assign n6709 = ~n6704 & n6708;
  assign n6710 = ~n6672 & n6709;
  assign n6711 = ~n6699 & ~n6707;
  assign n6712 = ~n6703 & ~n6711;
  assign n6713 = ~n6710 & ~n6712;
  assign n6714 = ~n6703 & n6708;
  assign n6715 = ~n6704 & n6714;
  assign n6716 = ~n6672 & ~n6711;
  assign n6717 = n6715 & n6716;
  assign n6718 = ~n6713 & ~n6717;
  assign n6719 = n6671 & ~n6718;
  assign n6720 = ~n6710 & n6712;
  assign n6721 = n6710 & ~n6712;
  assign n6722 = ~n6720 & ~n6721;
  assign n6723 = ~n6671 & ~n6722;
  assign n6724 = ~n6704 & ~n6707;
  assign n6725 = ~n6666 & ~n6672;
  assign n6726 = ~n6724 & n6725;
  assign n6727 = n6724 & ~n6725;
  assign n6728 = ~n6726 & ~n6727;
  assign n6729 = ~n6615 & ~n6618;
  assign n6730 = ~n6577 & ~n6583;
  assign n6731 = ~n6729 & n6730;
  assign n6732 = n6729 & ~n6730;
  assign n6733 = ~n6731 & ~n6732;
  assign n6734 = ~n6728 & ~n6733;
  assign n6735 = ~n6723 & ~n6734;
  assign n6736 = ~n6719 & n6735;
  assign n6737 = ~n6719 & ~n6723;
  assign n6738 = n6734 & ~n6737;
  assign n6739 = ~n6736 & ~n6738;
  assign n6740 = ~n6635 & ~n6739;
  assign n6741 = ~n6723 & n6734;
  assign n6742 = ~n6719 & n6741;
  assign n6743 = ~n6734 & ~n6737;
  assign n6744 = ~n6742 & ~n6743;
  assign n6745 = n6635 & ~n6744;
  assign n6746 = ~n6728 & n6733;
  assign n6747 = n6728 & ~n6733;
  assign n6748 = ~n6746 & ~n6747;
  assign n6749 = ~A193  & A194 ;
  assign n6750 = A193  & ~A194 ;
  assign n6751 = A195  & ~n6750;
  assign n6752 = ~n6749 & n6751;
  assign n6753 = ~n6749 & ~n6750;
  assign n6754 = ~A195  & ~n6753;
  assign n6755 = ~n6752 & ~n6754;
  assign n6756 = ~A196  & A197 ;
  assign n6757 = A196  & ~A197 ;
  assign n6758 = A198  & ~n6757;
  assign n6759 = ~n6756 & n6758;
  assign n6760 = ~n6756 & ~n6757;
  assign n6761 = ~A198  & ~n6760;
  assign n6762 = ~n6759 & ~n6761;
  assign n6763 = ~n6755 & n6762;
  assign n6764 = n6755 & ~n6762;
  assign n6765 = ~n6763 & ~n6764;
  assign n6766 = A196  & A197 ;
  assign n6767 = A198  & ~n6760;
  assign n6768 = ~n6766 & ~n6767;
  assign n6769 = A193  & A194 ;
  assign n6770 = A195  & ~n6753;
  assign n6771 = ~n6769 & ~n6770;
  assign n6772 = ~n6768 & n6771;
  assign n6773 = n6768 & ~n6771;
  assign n6774 = ~n6772 & ~n6773;
  assign n6775 = ~n6755 & ~n6762;
  assign n6776 = ~n6774 & n6775;
  assign n6777 = ~n6768 & ~n6771;
  assign n6778 = ~n6776 & ~n6777;
  assign n6779 = ~n6772 & n6775;
  assign n6780 = ~n6773 & n6779;
  assign n6781 = ~n6774 & ~n6775;
  assign n6782 = ~n6780 & ~n6781;
  assign n6783 = ~n6778 & ~n6782;
  assign n6784 = ~n6765 & ~n6783;
  assign n6785 = ~A187  & A188 ;
  assign n6786 = A187  & ~A188 ;
  assign n6787 = A189  & ~n6786;
  assign n6788 = ~n6785 & n6787;
  assign n6789 = ~n6785 & ~n6786;
  assign n6790 = ~A189  & ~n6789;
  assign n6791 = ~n6788 & ~n6790;
  assign n6792 = ~A190  & A191 ;
  assign n6793 = A190  & ~A191 ;
  assign n6794 = A192  & ~n6793;
  assign n6795 = ~n6792 & n6794;
  assign n6796 = ~n6792 & ~n6793;
  assign n6797 = ~A192  & ~n6796;
  assign n6798 = ~n6795 & ~n6797;
  assign n6799 = ~n6791 & n6798;
  assign n6800 = n6791 & ~n6798;
  assign n6801 = ~n6799 & ~n6800;
  assign n6802 = A190  & A191 ;
  assign n6803 = A192  & ~n6796;
  assign n6804 = ~n6802 & ~n6803;
  assign n6805 = A187  & A188 ;
  assign n6806 = A189  & ~n6789;
  assign n6807 = ~n6805 & ~n6806;
  assign n6808 = ~n6804 & n6807;
  assign n6809 = n6804 & ~n6807;
  assign n6810 = ~n6808 & ~n6809;
  assign n6811 = ~n6791 & ~n6798;
  assign n6812 = ~n6810 & n6811;
  assign n6813 = ~n6804 & ~n6807;
  assign n6814 = ~n6812 & ~n6813;
  assign n6815 = ~n6808 & n6811;
  assign n6816 = ~n6809 & n6815;
  assign n6817 = ~n6810 & ~n6811;
  assign n6818 = ~n6816 & ~n6817;
  assign n6819 = ~n6814 & ~n6818;
  assign n6820 = ~n6801 & ~n6819;
  assign n6821 = ~n6784 & n6820;
  assign n6822 = n6784 & ~n6820;
  assign n6823 = ~n6821 & ~n6822;
  assign n6824 = ~A181  & A182 ;
  assign n6825 = A181  & ~A182 ;
  assign n6826 = A183  & ~n6825;
  assign n6827 = ~n6824 & n6826;
  assign n6828 = ~n6824 & ~n6825;
  assign n6829 = ~A183  & ~n6828;
  assign n6830 = ~n6827 & ~n6829;
  assign n6831 = ~A184  & A185 ;
  assign n6832 = A184  & ~A185 ;
  assign n6833 = A186  & ~n6832;
  assign n6834 = ~n6831 & n6833;
  assign n6835 = ~n6831 & ~n6832;
  assign n6836 = ~A186  & ~n6835;
  assign n6837 = ~n6834 & ~n6836;
  assign n6838 = ~n6830 & n6837;
  assign n6839 = n6830 & ~n6837;
  assign n6840 = ~n6838 & ~n6839;
  assign n6841 = A184  & A185 ;
  assign n6842 = A186  & ~n6835;
  assign n6843 = ~n6841 & ~n6842;
  assign n6844 = A181  & A182 ;
  assign n6845 = A183  & ~n6828;
  assign n6846 = ~n6844 & ~n6845;
  assign n6847 = ~n6843 & n6846;
  assign n6848 = n6843 & ~n6846;
  assign n6849 = ~n6847 & ~n6848;
  assign n6850 = ~n6830 & ~n6837;
  assign n6851 = ~n6849 & n6850;
  assign n6852 = ~n6843 & ~n6846;
  assign n6853 = ~n6851 & ~n6852;
  assign n6854 = ~n6847 & n6850;
  assign n6855 = ~n6848 & n6854;
  assign n6856 = ~n6849 & ~n6850;
  assign n6857 = ~n6855 & ~n6856;
  assign n6858 = ~n6853 & ~n6857;
  assign n6859 = ~n6840 & ~n6858;
  assign n6860 = ~A175  & A176 ;
  assign n6861 = A175  & ~A176 ;
  assign n6862 = A177  & ~n6861;
  assign n6863 = ~n6860 & n6862;
  assign n6864 = ~n6860 & ~n6861;
  assign n6865 = ~A177  & ~n6864;
  assign n6866 = ~n6863 & ~n6865;
  assign n6867 = ~A178  & A179 ;
  assign n6868 = A178  & ~A179 ;
  assign n6869 = A180  & ~n6868;
  assign n6870 = ~n6867 & n6869;
  assign n6871 = ~n6867 & ~n6868;
  assign n6872 = ~A180  & ~n6871;
  assign n6873 = ~n6870 & ~n6872;
  assign n6874 = ~n6866 & n6873;
  assign n6875 = n6866 & ~n6873;
  assign n6876 = ~n6874 & ~n6875;
  assign n6877 = A178  & A179 ;
  assign n6878 = A180  & ~n6871;
  assign n6879 = ~n6877 & ~n6878;
  assign n6880 = A175  & A176 ;
  assign n6881 = A177  & ~n6864;
  assign n6882 = ~n6880 & ~n6881;
  assign n6883 = ~n6879 & n6882;
  assign n6884 = n6879 & ~n6882;
  assign n6885 = ~n6883 & ~n6884;
  assign n6886 = ~n6866 & ~n6873;
  assign n6887 = ~n6885 & n6886;
  assign n6888 = ~n6879 & ~n6882;
  assign n6889 = ~n6887 & ~n6888;
  assign n6890 = ~n6883 & n6886;
  assign n6891 = ~n6884 & n6890;
  assign n6892 = ~n6885 & ~n6886;
  assign n6893 = ~n6891 & ~n6892;
  assign n6894 = ~n6889 & ~n6893;
  assign n6895 = ~n6876 & ~n6894;
  assign n6896 = ~n6859 & n6895;
  assign n6897 = n6859 & ~n6895;
  assign n6898 = ~n6896 & ~n6897;
  assign n6899 = ~n6823 & n6898;
  assign n6900 = n6823 & ~n6898;
  assign n6901 = ~n6899 & ~n6900;
  assign n6902 = ~n6748 & ~n6901;
  assign n6903 = ~n6745 & n6902;
  assign n6904 = ~n6740 & n6903;
  assign n6905 = ~n6740 & ~n6745;
  assign n6906 = ~n6902 & ~n6905;
  assign n6907 = ~n6904 & ~n6906;
  assign n6908 = ~n6801 & ~n6814;
  assign n6909 = ~n6818 & ~n6908;
  assign n6910 = ~n6765 & ~n6801;
  assign n6911 = ~n6783 & n6910;
  assign n6912 = ~n6819 & n6911;
  assign n6913 = ~n6765 & ~n6778;
  assign n6914 = ~n6782 & ~n6913;
  assign n6915 = ~n6912 & ~n6914;
  assign n6916 = ~n6782 & n6910;
  assign n6917 = ~n6783 & n6916;
  assign n6918 = ~n6819 & ~n6913;
  assign n6919 = n6917 & n6918;
  assign n6920 = ~n6915 & ~n6919;
  assign n6921 = n6909 & ~n6920;
  assign n6922 = ~n6912 & n6914;
  assign n6923 = n6912 & ~n6914;
  assign n6924 = ~n6922 & ~n6923;
  assign n6925 = ~n6909 & ~n6924;
  assign n6926 = ~n6823 & ~n6898;
  assign n6927 = ~n6925 & n6926;
  assign n6928 = ~n6921 & n6927;
  assign n6929 = ~n6921 & ~n6925;
  assign n6930 = ~n6926 & ~n6929;
  assign n6931 = ~n6928 & ~n6930;
  assign n6932 = ~n6876 & ~n6889;
  assign n6933 = ~n6893 & ~n6932;
  assign n6934 = ~n6840 & ~n6876;
  assign n6935 = ~n6858 & n6934;
  assign n6936 = ~n6894 & n6935;
  assign n6937 = ~n6840 & ~n6853;
  assign n6938 = ~n6857 & ~n6937;
  assign n6939 = ~n6936 & n6938;
  assign n6940 = n6936 & ~n6938;
  assign n6941 = ~n6939 & ~n6940;
  assign n6942 = ~n6933 & ~n6941;
  assign n6943 = ~n6936 & ~n6938;
  assign n6944 = ~n6857 & n6934;
  assign n6945 = ~n6858 & n6944;
  assign n6946 = ~n6894 & ~n6937;
  assign n6947 = n6945 & n6946;
  assign n6948 = ~n6943 & ~n6947;
  assign n6949 = n6933 & ~n6948;
  assign n6950 = ~n6942 & ~n6949;
  assign n6951 = ~n6931 & n6950;
  assign n6952 = ~n6925 & ~n6926;
  assign n6953 = ~n6921 & n6952;
  assign n6954 = n6926 & ~n6929;
  assign n6955 = ~n6953 & ~n6954;
  assign n6956 = ~n6950 & ~n6955;
  assign n6957 = ~n6951 & ~n6956;
  assign n6958 = ~n6907 & n6957;
  assign n6959 = ~n6745 & ~n6902;
  assign n6960 = ~n6740 & n6959;
  assign n6961 = n6902 & ~n6905;
  assign n6962 = ~n6960 & ~n6961;
  assign n6963 = ~n6957 & ~n6962;
  assign n6964 = ~n6958 & ~n6963;
  assign n6965 = A238  & A239 ;
  assign n6966 = A238  & ~A239 ;
  assign n6967 = ~A238  & A239 ;
  assign n6968 = ~n6966 & ~n6967;
  assign n6969 = A240  & ~n6968;
  assign n6970 = ~n6965 & ~n6969;
  assign n6971 = A235  & A236 ;
  assign n6972 = A235  & ~A236 ;
  assign n6973 = ~A235  & A236 ;
  assign n6974 = ~n6972 & ~n6973;
  assign n6975 = A237  & ~n6974;
  assign n6976 = ~n6971 & ~n6975;
  assign n6977 = n6970 & ~n6976;
  assign n6978 = ~n6970 & n6976;
  assign n6979 = A237  & ~n6972;
  assign n6980 = ~n6973 & n6979;
  assign n6981 = ~A237  & ~n6974;
  assign n6982 = ~n6980 & ~n6981;
  assign n6983 = A240  & ~n6966;
  assign n6984 = ~n6967 & n6983;
  assign n6985 = ~A240  & ~n6968;
  assign n6986 = ~n6984 & ~n6985;
  assign n6987 = ~n6982 & ~n6986;
  assign n6988 = ~n6978 & n6987;
  assign n6989 = ~n6977 & n6988;
  assign n6990 = ~n6977 & ~n6978;
  assign n6991 = ~n6987 & ~n6990;
  assign n6992 = ~n6989 & ~n6991;
  assign n6993 = ~n6982 & n6986;
  assign n6994 = n6982 & ~n6986;
  assign n6995 = ~n6993 & ~n6994;
  assign n6996 = n6987 & ~n6990;
  assign n6997 = ~n6970 & ~n6976;
  assign n6998 = ~n6996 & ~n6997;
  assign n6999 = ~n6995 & ~n6998;
  assign n7000 = ~n6992 & ~n6999;
  assign n7001 = ~n6992 & ~n6998;
  assign n7002 = A244  & A245 ;
  assign n7003 = A244  & ~A245 ;
  assign n7004 = ~A244  & A245 ;
  assign n7005 = ~n7003 & ~n7004;
  assign n7006 = A246  & ~n7005;
  assign n7007 = ~n7002 & ~n7006;
  assign n7008 = A241  & A242 ;
  assign n7009 = A241  & ~A242 ;
  assign n7010 = ~A241  & A242 ;
  assign n7011 = ~n7009 & ~n7010;
  assign n7012 = A243  & ~n7011;
  assign n7013 = ~n7008 & ~n7012;
  assign n7014 = ~n7007 & n7013;
  assign n7015 = n7007 & ~n7013;
  assign n7016 = ~n7014 & ~n7015;
  assign n7017 = A243  & ~n7009;
  assign n7018 = ~n7010 & n7017;
  assign n7019 = ~A243  & ~n7011;
  assign n7020 = ~n7018 & ~n7019;
  assign n7021 = A246  & ~n7003;
  assign n7022 = ~n7004 & n7021;
  assign n7023 = ~A246  & ~n7005;
  assign n7024 = ~n7022 & ~n7023;
  assign n7025 = ~n7020 & ~n7024;
  assign n7026 = ~n7016 & n7025;
  assign n7027 = ~n7007 & ~n7013;
  assign n7028 = ~n7026 & ~n7027;
  assign n7029 = ~n7014 & n7025;
  assign n7030 = ~n7015 & n7029;
  assign n7031 = ~n7016 & ~n7025;
  assign n7032 = ~n7030 & ~n7031;
  assign n7033 = ~n7028 & ~n7032;
  assign n7034 = ~n7020 & n7024;
  assign n7035 = n7020 & ~n7024;
  assign n7036 = ~n7034 & ~n7035;
  assign n7037 = ~n6995 & ~n7036;
  assign n7038 = ~n7033 & n7037;
  assign n7039 = ~n7001 & n7038;
  assign n7040 = ~n7028 & ~n7036;
  assign n7041 = ~n7032 & ~n7040;
  assign n7042 = ~n7039 & ~n7041;
  assign n7043 = ~n7032 & n7037;
  assign n7044 = ~n7033 & n7043;
  assign n7045 = ~n7001 & ~n7040;
  assign n7046 = n7044 & n7045;
  assign n7047 = ~n7042 & ~n7046;
  assign n7048 = n7000 & ~n7047;
  assign n7049 = ~n7039 & n7041;
  assign n7050 = n7039 & ~n7041;
  assign n7051 = ~n7049 & ~n7050;
  assign n7052 = ~n7000 & ~n7051;
  assign n7053 = ~n7033 & ~n7036;
  assign n7054 = ~n6995 & ~n7001;
  assign n7055 = ~n7053 & n7054;
  assign n7056 = n7053 & ~n7054;
  assign n7057 = ~n7055 & ~n7056;
  assign n7058 = ~A229  & A230 ;
  assign n7059 = A229  & ~A230 ;
  assign n7060 = A231  & ~n7059;
  assign n7061 = ~n7058 & n7060;
  assign n7062 = ~n7058 & ~n7059;
  assign n7063 = ~A231  & ~n7062;
  assign n7064 = ~n7061 & ~n7063;
  assign n7065 = ~A232  & A233 ;
  assign n7066 = A232  & ~A233 ;
  assign n7067 = A234  & ~n7066;
  assign n7068 = ~n7065 & n7067;
  assign n7069 = ~n7065 & ~n7066;
  assign n7070 = ~A234  & ~n7069;
  assign n7071 = ~n7068 & ~n7070;
  assign n7072 = ~n7064 & n7071;
  assign n7073 = n7064 & ~n7071;
  assign n7074 = ~n7072 & ~n7073;
  assign n7075 = A232  & A233 ;
  assign n7076 = A234  & ~n7069;
  assign n7077 = ~n7075 & ~n7076;
  assign n7078 = A229  & A230 ;
  assign n7079 = A231  & ~n7062;
  assign n7080 = ~n7078 & ~n7079;
  assign n7081 = ~n7077 & n7080;
  assign n7082 = n7077 & ~n7080;
  assign n7083 = ~n7081 & ~n7082;
  assign n7084 = ~n7064 & ~n7071;
  assign n7085 = ~n7083 & n7084;
  assign n7086 = ~n7077 & ~n7080;
  assign n7087 = ~n7085 & ~n7086;
  assign n7088 = ~n7081 & n7084;
  assign n7089 = ~n7082 & n7088;
  assign n7090 = ~n7083 & ~n7084;
  assign n7091 = ~n7089 & ~n7090;
  assign n7092 = ~n7087 & ~n7091;
  assign n7093 = ~n7074 & ~n7092;
  assign n7094 = ~A223  & A224 ;
  assign n7095 = A223  & ~A224 ;
  assign n7096 = A225  & ~n7095;
  assign n7097 = ~n7094 & n7096;
  assign n7098 = ~n7094 & ~n7095;
  assign n7099 = ~A225  & ~n7098;
  assign n7100 = ~n7097 & ~n7099;
  assign n7101 = ~A226  & A227 ;
  assign n7102 = A226  & ~A227 ;
  assign n7103 = A228  & ~n7102;
  assign n7104 = ~n7101 & n7103;
  assign n7105 = ~n7101 & ~n7102;
  assign n7106 = ~A228  & ~n7105;
  assign n7107 = ~n7104 & ~n7106;
  assign n7108 = ~n7100 & n7107;
  assign n7109 = n7100 & ~n7107;
  assign n7110 = ~n7108 & ~n7109;
  assign n7111 = A226  & A227 ;
  assign n7112 = A228  & ~n7105;
  assign n7113 = ~n7111 & ~n7112;
  assign n7114 = A223  & A224 ;
  assign n7115 = A225  & ~n7098;
  assign n7116 = ~n7114 & ~n7115;
  assign n7117 = ~n7113 & n7116;
  assign n7118 = n7113 & ~n7116;
  assign n7119 = ~n7117 & ~n7118;
  assign n7120 = ~n7100 & ~n7107;
  assign n7121 = ~n7119 & n7120;
  assign n7122 = ~n7113 & ~n7116;
  assign n7123 = ~n7121 & ~n7122;
  assign n7124 = ~n7117 & n7120;
  assign n7125 = ~n7118 & n7124;
  assign n7126 = ~n7119 & ~n7120;
  assign n7127 = ~n7125 & ~n7126;
  assign n7128 = ~n7123 & ~n7127;
  assign n7129 = ~n7110 & ~n7128;
  assign n7130 = ~n7093 & n7129;
  assign n7131 = n7093 & ~n7129;
  assign n7132 = ~n7130 & ~n7131;
  assign n7133 = ~n7057 & ~n7132;
  assign n7134 = ~n7052 & n7133;
  assign n7135 = ~n7048 & n7134;
  assign n7136 = ~n7048 & ~n7052;
  assign n7137 = ~n7133 & ~n7136;
  assign n7138 = ~n7135 & ~n7137;
  assign n7139 = ~n7110 & ~n7123;
  assign n7140 = ~n7127 & ~n7139;
  assign n7141 = ~n7074 & ~n7110;
  assign n7142 = ~n7092 & n7141;
  assign n7143 = ~n7128 & n7142;
  assign n7144 = ~n7074 & ~n7087;
  assign n7145 = ~n7091 & ~n7144;
  assign n7146 = ~n7143 & n7145;
  assign n7147 = n7143 & ~n7145;
  assign n7148 = ~n7146 & ~n7147;
  assign n7149 = ~n7140 & ~n7148;
  assign n7150 = ~n7143 & ~n7145;
  assign n7151 = ~n7091 & n7141;
  assign n7152 = ~n7092 & n7151;
  assign n7153 = ~n7128 & ~n7144;
  assign n7154 = n7152 & n7153;
  assign n7155 = ~n7150 & ~n7154;
  assign n7156 = n7140 & ~n7155;
  assign n7157 = ~n7149 & ~n7156;
  assign n7158 = ~n7138 & n7157;
  assign n7159 = ~n7052 & ~n7133;
  assign n7160 = ~n7048 & n7159;
  assign n7161 = n7133 & ~n7136;
  assign n7162 = ~n7160 & ~n7161;
  assign n7163 = ~n7157 & ~n7162;
  assign n7164 = ~n7158 & ~n7163;
  assign n7165 = A250  & A251 ;
  assign n7166 = A250  & ~A251 ;
  assign n7167 = ~A250  & A251 ;
  assign n7168 = ~n7166 & ~n7167;
  assign n7169 = A252  & ~n7168;
  assign n7170 = ~n7165 & ~n7169;
  assign n7171 = A247  & A248 ;
  assign n7172 = A247  & ~A248 ;
  assign n7173 = ~A247  & A248 ;
  assign n7174 = ~n7172 & ~n7173;
  assign n7175 = A249  & ~n7174;
  assign n7176 = ~n7171 & ~n7175;
  assign n7177 = n7170 & ~n7176;
  assign n7178 = ~n7170 & n7176;
  assign n7179 = A249  & ~n7172;
  assign n7180 = ~n7173 & n7179;
  assign n7181 = ~A249  & ~n7174;
  assign n7182 = ~n7180 & ~n7181;
  assign n7183 = A252  & ~n7166;
  assign n7184 = ~n7167 & n7183;
  assign n7185 = ~A252  & ~n7168;
  assign n7186 = ~n7184 & ~n7185;
  assign n7187 = ~n7182 & ~n7186;
  assign n7188 = ~n7178 & n7187;
  assign n7189 = ~n7177 & n7188;
  assign n7190 = ~n7177 & ~n7178;
  assign n7191 = ~n7187 & ~n7190;
  assign n7192 = ~n7189 & ~n7191;
  assign n7193 = ~n7182 & n7186;
  assign n7194 = n7182 & ~n7186;
  assign n7195 = ~n7193 & ~n7194;
  assign n7196 = n7187 & ~n7190;
  assign n7197 = ~n7170 & ~n7176;
  assign n7198 = ~n7196 & ~n7197;
  assign n7199 = ~n7195 & ~n7198;
  assign n7200 = ~n7192 & ~n7199;
  assign n7201 = ~n7192 & ~n7198;
  assign n7202 = A256  & A257 ;
  assign n7203 = A256  & ~A257 ;
  assign n7204 = ~A256  & A257 ;
  assign n7205 = ~n7203 & ~n7204;
  assign n7206 = A258  & ~n7205;
  assign n7207 = ~n7202 & ~n7206;
  assign n7208 = A253  & A254 ;
  assign n7209 = A253  & ~A254 ;
  assign n7210 = ~A253  & A254 ;
  assign n7211 = ~n7209 & ~n7210;
  assign n7212 = A255  & ~n7211;
  assign n7213 = ~n7208 & ~n7212;
  assign n7214 = ~n7207 & n7213;
  assign n7215 = n7207 & ~n7213;
  assign n7216 = ~n7214 & ~n7215;
  assign n7217 = A255  & ~n7209;
  assign n7218 = ~n7210 & n7217;
  assign n7219 = ~A255  & ~n7211;
  assign n7220 = ~n7218 & ~n7219;
  assign n7221 = A258  & ~n7203;
  assign n7222 = ~n7204 & n7221;
  assign n7223 = ~A258  & ~n7205;
  assign n7224 = ~n7222 & ~n7223;
  assign n7225 = ~n7220 & ~n7224;
  assign n7226 = ~n7216 & n7225;
  assign n7227 = ~n7207 & ~n7213;
  assign n7228 = ~n7226 & ~n7227;
  assign n7229 = ~n7214 & n7225;
  assign n7230 = ~n7215 & n7229;
  assign n7231 = ~n7216 & ~n7225;
  assign n7232 = ~n7230 & ~n7231;
  assign n7233 = ~n7228 & ~n7232;
  assign n7234 = ~n7220 & n7224;
  assign n7235 = n7220 & ~n7224;
  assign n7236 = ~n7234 & ~n7235;
  assign n7237 = ~n7195 & ~n7236;
  assign n7238 = ~n7233 & n7237;
  assign n7239 = ~n7201 & n7238;
  assign n7240 = ~n7228 & ~n7236;
  assign n7241 = ~n7232 & ~n7240;
  assign n7242 = ~n7239 & n7241;
  assign n7243 = n7239 & ~n7241;
  assign n7244 = ~n7242 & ~n7243;
  assign n7245 = ~n7200 & ~n7244;
  assign n7246 = ~n7239 & ~n7241;
  assign n7247 = ~n7232 & n7237;
  assign n7248 = ~n7233 & n7247;
  assign n7249 = ~n7201 & ~n7240;
  assign n7250 = n7248 & n7249;
  assign n7251 = ~n7246 & ~n7250;
  assign n7252 = n7200 & ~n7251;
  assign n7253 = ~n7245 & ~n7252;
  assign n7254 = A262  & A263 ;
  assign n7255 = A262  & ~A263 ;
  assign n7256 = ~A262  & A263 ;
  assign n7257 = ~n7255 & ~n7256;
  assign n7258 = A264  & ~n7257;
  assign n7259 = ~n7254 & ~n7258;
  assign n7260 = A259  & A260 ;
  assign n7261 = A259  & ~A260 ;
  assign n7262 = ~A259  & A260 ;
  assign n7263 = ~n7261 & ~n7262;
  assign n7264 = A261  & ~n7263;
  assign n7265 = ~n7260 & ~n7264;
  assign n7266 = n7259 & ~n7265;
  assign n7267 = ~n7259 & n7265;
  assign n7268 = A261  & ~n7261;
  assign n7269 = ~n7262 & n7268;
  assign n7270 = ~A261  & ~n7263;
  assign n7271 = ~n7269 & ~n7270;
  assign n7272 = A264  & ~n7255;
  assign n7273 = ~n7256 & n7272;
  assign n7274 = ~A264  & ~n7257;
  assign n7275 = ~n7273 & ~n7274;
  assign n7276 = ~n7271 & ~n7275;
  assign n7277 = ~n7267 & n7276;
  assign n7278 = ~n7266 & n7277;
  assign n7279 = ~n7266 & ~n7267;
  assign n7280 = ~n7276 & ~n7279;
  assign n7281 = ~n7278 & ~n7280;
  assign n7282 = ~n7271 & n7275;
  assign n7283 = n7271 & ~n7275;
  assign n7284 = ~n7282 & ~n7283;
  assign n7285 = n7276 & ~n7279;
  assign n7286 = ~n7259 & ~n7265;
  assign n7287 = ~n7285 & ~n7286;
  assign n7288 = ~n7284 & ~n7287;
  assign n7289 = ~n7281 & ~n7288;
  assign n7290 = ~n7281 & ~n7287;
  assign n7291 = A268  & A269 ;
  assign n7292 = A268  & ~A269 ;
  assign n7293 = ~A268  & A269 ;
  assign n7294 = ~n7292 & ~n7293;
  assign n7295 = A270  & ~n7294;
  assign n7296 = ~n7291 & ~n7295;
  assign n7297 = A265  & A266 ;
  assign n7298 = A265  & ~A266 ;
  assign n7299 = ~A265  & A266 ;
  assign n7300 = ~n7298 & ~n7299;
  assign n7301 = A267  & ~n7300;
  assign n7302 = ~n7297 & ~n7301;
  assign n7303 = ~n7296 & n7302;
  assign n7304 = n7296 & ~n7302;
  assign n7305 = ~n7303 & ~n7304;
  assign n7306 = A267  & ~n7298;
  assign n7307 = ~n7299 & n7306;
  assign n7308 = ~A267  & ~n7300;
  assign n7309 = ~n7307 & ~n7308;
  assign n7310 = A270  & ~n7292;
  assign n7311 = ~n7293 & n7310;
  assign n7312 = ~A270  & ~n7294;
  assign n7313 = ~n7311 & ~n7312;
  assign n7314 = ~n7309 & ~n7313;
  assign n7315 = ~n7305 & n7314;
  assign n7316 = ~n7296 & ~n7302;
  assign n7317 = ~n7315 & ~n7316;
  assign n7318 = ~n7303 & n7314;
  assign n7319 = ~n7304 & n7318;
  assign n7320 = ~n7305 & ~n7314;
  assign n7321 = ~n7319 & ~n7320;
  assign n7322 = ~n7317 & ~n7321;
  assign n7323 = ~n7309 & n7313;
  assign n7324 = n7309 & ~n7313;
  assign n7325 = ~n7323 & ~n7324;
  assign n7326 = ~n7284 & ~n7325;
  assign n7327 = ~n7322 & n7326;
  assign n7328 = ~n7290 & n7327;
  assign n7329 = ~n7317 & ~n7325;
  assign n7330 = ~n7321 & ~n7329;
  assign n7331 = ~n7328 & ~n7330;
  assign n7332 = ~n7321 & n7326;
  assign n7333 = ~n7322 & n7332;
  assign n7334 = ~n7290 & ~n7329;
  assign n7335 = n7333 & n7334;
  assign n7336 = ~n7331 & ~n7335;
  assign n7337 = n7289 & ~n7336;
  assign n7338 = ~n7328 & n7330;
  assign n7339 = n7328 & ~n7330;
  assign n7340 = ~n7338 & ~n7339;
  assign n7341 = ~n7289 & ~n7340;
  assign n7342 = ~n7322 & ~n7325;
  assign n7343 = ~n7284 & ~n7290;
  assign n7344 = ~n7342 & n7343;
  assign n7345 = n7342 & ~n7343;
  assign n7346 = ~n7344 & ~n7345;
  assign n7347 = ~n7233 & ~n7236;
  assign n7348 = ~n7195 & ~n7201;
  assign n7349 = ~n7347 & n7348;
  assign n7350 = n7347 & ~n7348;
  assign n7351 = ~n7349 & ~n7350;
  assign n7352 = ~n7346 & ~n7351;
  assign n7353 = ~n7341 & ~n7352;
  assign n7354 = ~n7337 & n7353;
  assign n7355 = ~n7337 & ~n7341;
  assign n7356 = n7352 & ~n7355;
  assign n7357 = ~n7354 & ~n7356;
  assign n7358 = ~n7253 & ~n7357;
  assign n7359 = ~n7341 & n7352;
  assign n7360 = ~n7337 & n7359;
  assign n7361 = ~n7352 & ~n7355;
  assign n7362 = ~n7360 & ~n7361;
  assign n7363 = n7253 & ~n7362;
  assign n7364 = ~n7346 & n7351;
  assign n7365 = n7346 & ~n7351;
  assign n7366 = ~n7364 & ~n7365;
  assign n7367 = ~n7057 & n7132;
  assign n7368 = n7057 & ~n7132;
  assign n7369 = ~n7367 & ~n7368;
  assign n7370 = ~n7366 & ~n7369;
  assign n7371 = ~n7363 & ~n7370;
  assign n7372 = ~n7358 & n7371;
  assign n7373 = ~n7358 & ~n7363;
  assign n7374 = n7370 & ~n7373;
  assign n7375 = ~n7372 & ~n7374;
  assign n7376 = ~n7164 & ~n7375;
  assign n7377 = ~n7363 & n7370;
  assign n7378 = ~n7358 & n7377;
  assign n7379 = ~n7370 & ~n7373;
  assign n7380 = ~n7378 & ~n7379;
  assign n7381 = n7164 & ~n7380;
  assign n7382 = ~n7366 & n7369;
  assign n7383 = n7366 & ~n7369;
  assign n7384 = ~n7382 & ~n7383;
  assign n7385 = ~n6748 & n6901;
  assign n7386 = n6748 & ~n6901;
  assign n7387 = ~n7385 & ~n7386;
  assign n7388 = ~n7384 & ~n7387;
  assign n7389 = ~n7381 & ~n7388;
  assign n7390 = ~n7376 & n7389;
  assign n7391 = ~n7376 & ~n7381;
  assign n7392 = n7388 & ~n7391;
  assign n7393 = ~n7390 & ~n7392;
  assign n7394 = ~n6964 & ~n7393;
  assign n7395 = ~n7381 & n7388;
  assign n7396 = ~n7376 & n7395;
  assign n7397 = ~n7388 & ~n7391;
  assign n7398 = ~n7396 & ~n7397;
  assign n7399 = n6964 & ~n7398;
  assign n7400 = ~n7384 & n7387;
  assign n7401 = n7384 & ~n7387;
  assign n7402 = ~n7400 & ~n7401;
  assign n7403 = ~A169  & A170 ;
  assign n7404 = A169  & ~A170 ;
  assign n7405 = A171  & ~n7404;
  assign n7406 = ~n7403 & n7405;
  assign n7407 = ~n7403 & ~n7404;
  assign n7408 = ~A171  & ~n7407;
  assign n7409 = ~n7406 & ~n7408;
  assign n7410 = ~A172  & A173 ;
  assign n7411 = A172  & ~A173 ;
  assign n7412 = A174  & ~n7411;
  assign n7413 = ~n7410 & n7412;
  assign n7414 = ~n7410 & ~n7411;
  assign n7415 = ~A174  & ~n7414;
  assign n7416 = ~n7413 & ~n7415;
  assign n7417 = ~n7409 & n7416;
  assign n7418 = n7409 & ~n7416;
  assign n7419 = ~n7417 & ~n7418;
  assign n7420 = A172  & A173 ;
  assign n7421 = A174  & ~n7414;
  assign n7422 = ~n7420 & ~n7421;
  assign n7423 = A169  & A170 ;
  assign n7424 = A171  & ~n7407;
  assign n7425 = ~n7423 & ~n7424;
  assign n7426 = ~n7422 & n7425;
  assign n7427 = n7422 & ~n7425;
  assign n7428 = ~n7426 & ~n7427;
  assign n7429 = ~n7409 & ~n7416;
  assign n7430 = ~n7428 & n7429;
  assign n7431 = ~n7422 & ~n7425;
  assign n7432 = ~n7430 & ~n7431;
  assign n7433 = ~n7426 & n7429;
  assign n7434 = ~n7427 & n7433;
  assign n7435 = ~n7428 & ~n7429;
  assign n7436 = ~n7434 & ~n7435;
  assign n7437 = ~n7432 & ~n7436;
  assign n7438 = ~n7419 & ~n7437;
  assign n7439 = ~A163  & A164 ;
  assign n7440 = A163  & ~A164 ;
  assign n7441 = A165  & ~n7440;
  assign n7442 = ~n7439 & n7441;
  assign n7443 = ~n7439 & ~n7440;
  assign n7444 = ~A165  & ~n7443;
  assign n7445 = ~n7442 & ~n7444;
  assign n7446 = ~A166  & A167 ;
  assign n7447 = A166  & ~A167 ;
  assign n7448 = A168  & ~n7447;
  assign n7449 = ~n7446 & n7448;
  assign n7450 = ~n7446 & ~n7447;
  assign n7451 = ~A168  & ~n7450;
  assign n7452 = ~n7449 & ~n7451;
  assign n7453 = ~n7445 & n7452;
  assign n7454 = n7445 & ~n7452;
  assign n7455 = ~n7453 & ~n7454;
  assign n7456 = A166  & A167 ;
  assign n7457 = A168  & ~n7450;
  assign n7458 = ~n7456 & ~n7457;
  assign n7459 = A163  & A164 ;
  assign n7460 = A165  & ~n7443;
  assign n7461 = ~n7459 & ~n7460;
  assign n7462 = ~n7458 & n7461;
  assign n7463 = n7458 & ~n7461;
  assign n7464 = ~n7462 & ~n7463;
  assign n7465 = ~n7445 & ~n7452;
  assign n7466 = ~n7464 & n7465;
  assign n7467 = ~n7458 & ~n7461;
  assign n7468 = ~n7466 & ~n7467;
  assign n7469 = ~n7462 & n7465;
  assign n7470 = ~n7463 & n7469;
  assign n7471 = ~n7464 & ~n7465;
  assign n7472 = ~n7470 & ~n7471;
  assign n7473 = ~n7468 & ~n7472;
  assign n7474 = ~n7455 & ~n7473;
  assign n7475 = ~n7438 & n7474;
  assign n7476 = n7438 & ~n7474;
  assign n7477 = ~n7475 & ~n7476;
  assign n7478 = ~A157  & A158 ;
  assign n7479 = A157  & ~A158 ;
  assign n7480 = A159  & ~n7479;
  assign n7481 = ~n7478 & n7480;
  assign n7482 = ~n7478 & ~n7479;
  assign n7483 = ~A159  & ~n7482;
  assign n7484 = ~n7481 & ~n7483;
  assign n7485 = ~A160  & A161 ;
  assign n7486 = A160  & ~A161 ;
  assign n7487 = A162  & ~n7486;
  assign n7488 = ~n7485 & n7487;
  assign n7489 = ~n7485 & ~n7486;
  assign n7490 = ~A162  & ~n7489;
  assign n7491 = ~n7488 & ~n7490;
  assign n7492 = ~n7484 & n7491;
  assign n7493 = n7484 & ~n7491;
  assign n7494 = ~n7492 & ~n7493;
  assign n7495 = A160  & A161 ;
  assign n7496 = A162  & ~n7489;
  assign n7497 = ~n7495 & ~n7496;
  assign n7498 = A157  & A158 ;
  assign n7499 = A159  & ~n7482;
  assign n7500 = ~n7498 & ~n7499;
  assign n7501 = ~n7497 & n7500;
  assign n7502 = n7497 & ~n7500;
  assign n7503 = ~n7501 & ~n7502;
  assign n7504 = ~n7484 & ~n7491;
  assign n7505 = ~n7503 & n7504;
  assign n7506 = ~n7497 & ~n7500;
  assign n7507 = ~n7505 & ~n7506;
  assign n7508 = ~n7501 & n7504;
  assign n7509 = ~n7502 & n7508;
  assign n7510 = ~n7503 & ~n7504;
  assign n7511 = ~n7509 & ~n7510;
  assign n7512 = ~n7507 & ~n7511;
  assign n7513 = ~n7494 & ~n7512;
  assign n7514 = ~A151  & A152 ;
  assign n7515 = A151  & ~A152 ;
  assign n7516 = A153  & ~n7515;
  assign n7517 = ~n7514 & n7516;
  assign n7518 = ~n7514 & ~n7515;
  assign n7519 = ~A153  & ~n7518;
  assign n7520 = ~n7517 & ~n7519;
  assign n7521 = ~A154  & A155 ;
  assign n7522 = A154  & ~A155 ;
  assign n7523 = A156  & ~n7522;
  assign n7524 = ~n7521 & n7523;
  assign n7525 = ~n7521 & ~n7522;
  assign n7526 = ~A156  & ~n7525;
  assign n7527 = ~n7524 & ~n7526;
  assign n7528 = ~n7520 & n7527;
  assign n7529 = n7520 & ~n7527;
  assign n7530 = ~n7528 & ~n7529;
  assign n7531 = A154  & A155 ;
  assign n7532 = A156  & ~n7525;
  assign n7533 = ~n7531 & ~n7532;
  assign n7534 = A151  & A152 ;
  assign n7535 = A153  & ~n7518;
  assign n7536 = ~n7534 & ~n7535;
  assign n7537 = ~n7533 & n7536;
  assign n7538 = n7533 & ~n7536;
  assign n7539 = ~n7537 & ~n7538;
  assign n7540 = ~n7520 & ~n7527;
  assign n7541 = ~n7539 & n7540;
  assign n7542 = ~n7533 & ~n7536;
  assign n7543 = ~n7541 & ~n7542;
  assign n7544 = ~n7537 & n7540;
  assign n7545 = ~n7538 & n7544;
  assign n7546 = ~n7539 & ~n7540;
  assign n7547 = ~n7545 & ~n7546;
  assign n7548 = ~n7543 & ~n7547;
  assign n7549 = ~n7530 & ~n7548;
  assign n7550 = ~n7513 & n7549;
  assign n7551 = n7513 & ~n7549;
  assign n7552 = ~n7550 & ~n7551;
  assign n7553 = ~n7477 & n7552;
  assign n7554 = n7477 & ~n7552;
  assign n7555 = ~n7553 & ~n7554;
  assign n7556 = ~A145  & A146 ;
  assign n7557 = A145  & ~A146 ;
  assign n7558 = A147  & ~n7557;
  assign n7559 = ~n7556 & n7558;
  assign n7560 = ~n7556 & ~n7557;
  assign n7561 = ~A147  & ~n7560;
  assign n7562 = ~n7559 & ~n7561;
  assign n7563 = ~A148  & A149 ;
  assign n7564 = A148  & ~A149 ;
  assign n7565 = A150  & ~n7564;
  assign n7566 = ~n7563 & n7565;
  assign n7567 = ~n7563 & ~n7564;
  assign n7568 = ~A150  & ~n7567;
  assign n7569 = ~n7566 & ~n7568;
  assign n7570 = ~n7562 & n7569;
  assign n7571 = n7562 & ~n7569;
  assign n7572 = ~n7570 & ~n7571;
  assign n7573 = A148  & A149 ;
  assign n7574 = A150  & ~n7567;
  assign n7575 = ~n7573 & ~n7574;
  assign n7576 = A145  & A146 ;
  assign n7577 = A147  & ~n7560;
  assign n7578 = ~n7576 & ~n7577;
  assign n7579 = ~n7575 & n7578;
  assign n7580 = n7575 & ~n7578;
  assign n7581 = ~n7579 & ~n7580;
  assign n7582 = ~n7562 & ~n7569;
  assign n7583 = ~n7581 & n7582;
  assign n7584 = ~n7575 & ~n7578;
  assign n7585 = ~n7583 & ~n7584;
  assign n7586 = ~n7579 & n7582;
  assign n7587 = ~n7580 & n7586;
  assign n7588 = ~n7581 & ~n7582;
  assign n7589 = ~n7587 & ~n7588;
  assign n7590 = ~n7585 & ~n7589;
  assign n7591 = ~n7572 & ~n7590;
  assign n7592 = ~A139  & A140 ;
  assign n7593 = A139  & ~A140 ;
  assign n7594 = A141  & ~n7593;
  assign n7595 = ~n7592 & n7594;
  assign n7596 = ~n7592 & ~n7593;
  assign n7597 = ~A141  & ~n7596;
  assign n7598 = ~n7595 & ~n7597;
  assign n7599 = ~A142  & A143 ;
  assign n7600 = A142  & ~A143 ;
  assign n7601 = A144  & ~n7600;
  assign n7602 = ~n7599 & n7601;
  assign n7603 = ~n7599 & ~n7600;
  assign n7604 = ~A144  & ~n7603;
  assign n7605 = ~n7602 & ~n7604;
  assign n7606 = ~n7598 & n7605;
  assign n7607 = n7598 & ~n7605;
  assign n7608 = ~n7606 & ~n7607;
  assign n7609 = A142  & A143 ;
  assign n7610 = A144  & ~n7603;
  assign n7611 = ~n7609 & ~n7610;
  assign n7612 = A139  & A140 ;
  assign n7613 = A141  & ~n7596;
  assign n7614 = ~n7612 & ~n7613;
  assign n7615 = ~n7611 & n7614;
  assign n7616 = n7611 & ~n7614;
  assign n7617 = ~n7615 & ~n7616;
  assign n7618 = ~n7598 & ~n7605;
  assign n7619 = ~n7617 & n7618;
  assign n7620 = ~n7611 & ~n7614;
  assign n7621 = ~n7619 & ~n7620;
  assign n7622 = ~n7615 & n7618;
  assign n7623 = ~n7616 & n7622;
  assign n7624 = ~n7617 & ~n7618;
  assign n7625 = ~n7623 & ~n7624;
  assign n7626 = ~n7621 & ~n7625;
  assign n7627 = ~n7608 & ~n7626;
  assign n7628 = ~n7591 & n7627;
  assign n7629 = n7591 & ~n7627;
  assign n7630 = ~n7628 & ~n7629;
  assign n7631 = ~A133  & A134 ;
  assign n7632 = A133  & ~A134 ;
  assign n7633 = A135  & ~n7632;
  assign n7634 = ~n7631 & n7633;
  assign n7635 = ~n7631 & ~n7632;
  assign n7636 = ~A135  & ~n7635;
  assign n7637 = ~n7634 & ~n7636;
  assign n7638 = ~A136  & A137 ;
  assign n7639 = A136  & ~A137 ;
  assign n7640 = A138  & ~n7639;
  assign n7641 = ~n7638 & n7640;
  assign n7642 = ~n7638 & ~n7639;
  assign n7643 = ~A138  & ~n7642;
  assign n7644 = ~n7641 & ~n7643;
  assign n7645 = ~n7637 & n7644;
  assign n7646 = n7637 & ~n7644;
  assign n7647 = ~n7645 & ~n7646;
  assign n7648 = A136  & A137 ;
  assign n7649 = A138  & ~n7642;
  assign n7650 = ~n7648 & ~n7649;
  assign n7651 = A133  & A134 ;
  assign n7652 = A135  & ~n7635;
  assign n7653 = ~n7651 & ~n7652;
  assign n7654 = ~n7650 & n7653;
  assign n7655 = n7650 & ~n7653;
  assign n7656 = ~n7654 & ~n7655;
  assign n7657 = ~n7637 & ~n7644;
  assign n7658 = ~n7656 & n7657;
  assign n7659 = ~n7650 & ~n7653;
  assign n7660 = ~n7658 & ~n7659;
  assign n7661 = ~n7654 & n7657;
  assign n7662 = ~n7655 & n7661;
  assign n7663 = ~n7656 & ~n7657;
  assign n7664 = ~n7662 & ~n7663;
  assign n7665 = ~n7660 & ~n7664;
  assign n7666 = ~n7647 & ~n7665;
  assign n7667 = ~A127  & A128 ;
  assign n7668 = A127  & ~A128 ;
  assign n7669 = A129  & ~n7668;
  assign n7670 = ~n7667 & n7669;
  assign n7671 = ~n7667 & ~n7668;
  assign n7672 = ~A129  & ~n7671;
  assign n7673 = ~n7670 & ~n7672;
  assign n7674 = ~A130  & A131 ;
  assign n7675 = A130  & ~A131 ;
  assign n7676 = A132  & ~n7675;
  assign n7677 = ~n7674 & n7676;
  assign n7678 = ~n7674 & ~n7675;
  assign n7679 = ~A132  & ~n7678;
  assign n7680 = ~n7677 & ~n7679;
  assign n7681 = ~n7673 & n7680;
  assign n7682 = n7673 & ~n7680;
  assign n7683 = ~n7681 & ~n7682;
  assign n7684 = A130  & A131 ;
  assign n7685 = A132  & ~n7678;
  assign n7686 = ~n7684 & ~n7685;
  assign n7687 = A127  & A128 ;
  assign n7688 = A129  & ~n7671;
  assign n7689 = ~n7687 & ~n7688;
  assign n7690 = ~n7686 & n7689;
  assign n7691 = n7686 & ~n7689;
  assign n7692 = ~n7690 & ~n7691;
  assign n7693 = ~n7673 & ~n7680;
  assign n7694 = ~n7692 & n7693;
  assign n7695 = ~n7686 & ~n7689;
  assign n7696 = ~n7694 & ~n7695;
  assign n7697 = ~n7690 & n7693;
  assign n7698 = ~n7691 & n7697;
  assign n7699 = ~n7692 & ~n7693;
  assign n7700 = ~n7698 & ~n7699;
  assign n7701 = ~n7696 & ~n7700;
  assign n7702 = ~n7683 & ~n7701;
  assign n7703 = ~n7666 & n7702;
  assign n7704 = n7666 & ~n7702;
  assign n7705 = ~n7703 & ~n7704;
  assign n7706 = ~n7630 & n7705;
  assign n7707 = n7630 & ~n7705;
  assign n7708 = ~n7706 & ~n7707;
  assign n7709 = ~n7555 & n7708;
  assign n7710 = n7555 & ~n7708;
  assign n7711 = ~n7709 & ~n7710;
  assign n7712 = ~A121  & A122 ;
  assign n7713 = A121  & ~A122 ;
  assign n7714 = A123  & ~n7713;
  assign n7715 = ~n7712 & n7714;
  assign n7716 = ~n7712 & ~n7713;
  assign n7717 = ~A123  & ~n7716;
  assign n7718 = ~n7715 & ~n7717;
  assign n7719 = ~A124  & A125 ;
  assign n7720 = A124  & ~A125 ;
  assign n7721 = A126  & ~n7720;
  assign n7722 = ~n7719 & n7721;
  assign n7723 = ~n7719 & ~n7720;
  assign n7724 = ~A126  & ~n7723;
  assign n7725 = ~n7722 & ~n7724;
  assign n7726 = ~n7718 & n7725;
  assign n7727 = n7718 & ~n7725;
  assign n7728 = ~n7726 & ~n7727;
  assign n7729 = A124  & A125 ;
  assign n7730 = A126  & ~n7723;
  assign n7731 = ~n7729 & ~n7730;
  assign n7732 = A121  & A122 ;
  assign n7733 = A123  & ~n7716;
  assign n7734 = ~n7732 & ~n7733;
  assign n7735 = ~n7731 & n7734;
  assign n7736 = n7731 & ~n7734;
  assign n7737 = ~n7735 & ~n7736;
  assign n7738 = ~n7718 & ~n7725;
  assign n7739 = ~n7737 & n7738;
  assign n7740 = ~n7731 & ~n7734;
  assign n7741 = ~n7739 & ~n7740;
  assign n7742 = ~n7735 & n7738;
  assign n7743 = ~n7736 & n7742;
  assign n7744 = ~n7737 & ~n7738;
  assign n7745 = ~n7743 & ~n7744;
  assign n7746 = ~n7741 & ~n7745;
  assign n7747 = ~n7728 & ~n7746;
  assign n7748 = ~A115  & A116 ;
  assign n7749 = A115  & ~A116 ;
  assign n7750 = A117  & ~n7749;
  assign n7751 = ~n7748 & n7750;
  assign n7752 = ~n7748 & ~n7749;
  assign n7753 = ~A117  & ~n7752;
  assign n7754 = ~n7751 & ~n7753;
  assign n7755 = ~A118  & A119 ;
  assign n7756 = A118  & ~A119 ;
  assign n7757 = A120  & ~n7756;
  assign n7758 = ~n7755 & n7757;
  assign n7759 = ~n7755 & ~n7756;
  assign n7760 = ~A120  & ~n7759;
  assign n7761 = ~n7758 & ~n7760;
  assign n7762 = ~n7754 & n7761;
  assign n7763 = n7754 & ~n7761;
  assign n7764 = ~n7762 & ~n7763;
  assign n7765 = A118  & A119 ;
  assign n7766 = A120  & ~n7759;
  assign n7767 = ~n7765 & ~n7766;
  assign n7768 = A115  & A116 ;
  assign n7769 = A117  & ~n7752;
  assign n7770 = ~n7768 & ~n7769;
  assign n7771 = ~n7767 & n7770;
  assign n7772 = n7767 & ~n7770;
  assign n7773 = ~n7771 & ~n7772;
  assign n7774 = ~n7754 & ~n7761;
  assign n7775 = ~n7773 & n7774;
  assign n7776 = ~n7767 & ~n7770;
  assign n7777 = ~n7775 & ~n7776;
  assign n7778 = ~n7771 & n7774;
  assign n7779 = ~n7772 & n7778;
  assign n7780 = ~n7773 & ~n7774;
  assign n7781 = ~n7779 & ~n7780;
  assign n7782 = ~n7777 & ~n7781;
  assign n7783 = ~n7764 & ~n7782;
  assign n7784 = ~n7747 & n7783;
  assign n7785 = n7747 & ~n7783;
  assign n7786 = ~n7784 & ~n7785;
  assign n7787 = ~A109  & A110 ;
  assign n7788 = A109  & ~A110 ;
  assign n7789 = A111  & ~n7788;
  assign n7790 = ~n7787 & n7789;
  assign n7791 = ~n7787 & ~n7788;
  assign n7792 = ~A111  & ~n7791;
  assign n7793 = ~n7790 & ~n7792;
  assign n7794 = ~A112  & A113 ;
  assign n7795 = A112  & ~A113 ;
  assign n7796 = A114  & ~n7795;
  assign n7797 = ~n7794 & n7796;
  assign n7798 = ~n7794 & ~n7795;
  assign n7799 = ~A114  & ~n7798;
  assign n7800 = ~n7797 & ~n7799;
  assign n7801 = ~n7793 & n7800;
  assign n7802 = n7793 & ~n7800;
  assign n7803 = ~n7801 & ~n7802;
  assign n7804 = A112  & A113 ;
  assign n7805 = A114  & ~n7798;
  assign n7806 = ~n7804 & ~n7805;
  assign n7807 = A109  & A110 ;
  assign n7808 = A111  & ~n7791;
  assign n7809 = ~n7807 & ~n7808;
  assign n7810 = ~n7806 & n7809;
  assign n7811 = n7806 & ~n7809;
  assign n7812 = ~n7810 & ~n7811;
  assign n7813 = ~n7793 & ~n7800;
  assign n7814 = ~n7812 & n7813;
  assign n7815 = ~n7806 & ~n7809;
  assign n7816 = ~n7814 & ~n7815;
  assign n7817 = ~n7810 & n7813;
  assign n7818 = ~n7811 & n7817;
  assign n7819 = ~n7812 & ~n7813;
  assign n7820 = ~n7818 & ~n7819;
  assign n7821 = ~n7816 & ~n7820;
  assign n7822 = ~n7803 & ~n7821;
  assign n7823 = ~A103  & A104 ;
  assign n7824 = A103  & ~A104 ;
  assign n7825 = A105  & ~n7824;
  assign n7826 = ~n7823 & n7825;
  assign n7827 = ~n7823 & ~n7824;
  assign n7828 = ~A105  & ~n7827;
  assign n7829 = ~n7826 & ~n7828;
  assign n7830 = ~A106  & A107 ;
  assign n7831 = A106  & ~A107 ;
  assign n7832 = A108  & ~n7831;
  assign n7833 = ~n7830 & n7832;
  assign n7834 = ~n7830 & ~n7831;
  assign n7835 = ~A108  & ~n7834;
  assign n7836 = ~n7833 & ~n7835;
  assign n7837 = ~n7829 & n7836;
  assign n7838 = n7829 & ~n7836;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = A106  & A107 ;
  assign n7841 = A108  & ~n7834;
  assign n7842 = ~n7840 & ~n7841;
  assign n7843 = A103  & A104 ;
  assign n7844 = A105  & ~n7827;
  assign n7845 = ~n7843 & ~n7844;
  assign n7846 = ~n7842 & n7845;
  assign n7847 = n7842 & ~n7845;
  assign n7848 = ~n7846 & ~n7847;
  assign n7849 = ~n7829 & ~n7836;
  assign n7850 = ~n7848 & n7849;
  assign n7851 = ~n7842 & ~n7845;
  assign n7852 = ~n7850 & ~n7851;
  assign n7853 = ~n7846 & n7849;
  assign n7854 = ~n7847 & n7853;
  assign n7855 = ~n7848 & ~n7849;
  assign n7856 = ~n7854 & ~n7855;
  assign n7857 = ~n7852 & ~n7856;
  assign n7858 = ~n7839 & ~n7857;
  assign n7859 = ~n7822 & n7858;
  assign n7860 = n7822 & ~n7858;
  assign n7861 = ~n7859 & ~n7860;
  assign n7862 = ~n7786 & n7861;
  assign n7863 = n7786 & ~n7861;
  assign n7864 = ~n7862 & ~n7863;
  assign n7865 = ~A97  & A98 ;
  assign n7866 = A97  & ~A98 ;
  assign n7867 = A99  & ~n7866;
  assign n7868 = ~n7865 & n7867;
  assign n7869 = ~n7865 & ~n7866;
  assign n7870 = ~A99  & ~n7869;
  assign n7871 = ~n7868 & ~n7870;
  assign n7872 = ~A100  & A101 ;
  assign n7873 = A100  & ~A101 ;
  assign n7874 = A102  & ~n7873;
  assign n7875 = ~n7872 & n7874;
  assign n7876 = ~n7872 & ~n7873;
  assign n7877 = ~A102  & ~n7876;
  assign n7878 = ~n7875 & ~n7877;
  assign n7879 = ~n7871 & n7878;
  assign n7880 = n7871 & ~n7878;
  assign n7881 = ~n7879 & ~n7880;
  assign n7882 = A100  & A101 ;
  assign n7883 = A102  & ~n7876;
  assign n7884 = ~n7882 & ~n7883;
  assign n7885 = A97  & A98 ;
  assign n7886 = A99  & ~n7869;
  assign n7887 = ~n7885 & ~n7886;
  assign n7888 = ~n7884 & n7887;
  assign n7889 = n7884 & ~n7887;
  assign n7890 = ~n7888 & ~n7889;
  assign n7891 = ~n7871 & ~n7878;
  assign n7892 = ~n7890 & n7891;
  assign n7893 = ~n7884 & ~n7887;
  assign n7894 = ~n7892 & ~n7893;
  assign n7895 = ~n7888 & n7891;
  assign n7896 = ~n7889 & n7895;
  assign n7897 = ~n7890 & ~n7891;
  assign n7898 = ~n7896 & ~n7897;
  assign n7899 = ~n7894 & ~n7898;
  assign n7900 = ~n7881 & ~n7899;
  assign n7901 = ~A91  & A92 ;
  assign n7902 = A91  & ~A92 ;
  assign n7903 = A93  & ~n7902;
  assign n7904 = ~n7901 & n7903;
  assign n7905 = ~n7901 & ~n7902;
  assign n7906 = ~A93  & ~n7905;
  assign n7907 = ~n7904 & ~n7906;
  assign n7908 = ~A94  & A95 ;
  assign n7909 = A94  & ~A95 ;
  assign n7910 = A96  & ~n7909;
  assign n7911 = ~n7908 & n7910;
  assign n7912 = ~n7908 & ~n7909;
  assign n7913 = ~A96  & ~n7912;
  assign n7914 = ~n7911 & ~n7913;
  assign n7915 = ~n7907 & n7914;
  assign n7916 = n7907 & ~n7914;
  assign n7917 = ~n7915 & ~n7916;
  assign n7918 = A94  & A95 ;
  assign n7919 = A96  & ~n7912;
  assign n7920 = ~n7918 & ~n7919;
  assign n7921 = A91  & A92 ;
  assign n7922 = A93  & ~n7905;
  assign n7923 = ~n7921 & ~n7922;
  assign n7924 = ~n7920 & n7923;
  assign n7925 = n7920 & ~n7923;
  assign n7926 = ~n7924 & ~n7925;
  assign n7927 = ~n7907 & ~n7914;
  assign n7928 = ~n7926 & n7927;
  assign n7929 = ~n7920 & ~n7923;
  assign n7930 = ~n7928 & ~n7929;
  assign n7931 = ~n7924 & n7927;
  assign n7932 = ~n7925 & n7931;
  assign n7933 = ~n7926 & ~n7927;
  assign n7934 = ~n7932 & ~n7933;
  assign n7935 = ~n7930 & ~n7934;
  assign n7936 = ~n7917 & ~n7935;
  assign n7937 = ~n7900 & n7936;
  assign n7938 = n7900 & ~n7936;
  assign n7939 = ~n7937 & ~n7938;
  assign n7940 = ~A85  & A86 ;
  assign n7941 = A85  & ~A86 ;
  assign n7942 = A87  & ~n7941;
  assign n7943 = ~n7940 & n7942;
  assign n7944 = ~n7940 & ~n7941;
  assign n7945 = ~A87  & ~n7944;
  assign n7946 = ~n7943 & ~n7945;
  assign n7947 = ~A88  & A89 ;
  assign n7948 = A88  & ~A89 ;
  assign n7949 = A90  & ~n7948;
  assign n7950 = ~n7947 & n7949;
  assign n7951 = ~n7947 & ~n7948;
  assign n7952 = ~A90  & ~n7951;
  assign n7953 = ~n7950 & ~n7952;
  assign n7954 = ~n7946 & n7953;
  assign n7955 = n7946 & ~n7953;
  assign n7956 = ~n7954 & ~n7955;
  assign n7957 = A88  & A89 ;
  assign n7958 = A90  & ~n7951;
  assign n7959 = ~n7957 & ~n7958;
  assign n7960 = A85  & A86 ;
  assign n7961 = A87  & ~n7944;
  assign n7962 = ~n7960 & ~n7961;
  assign n7963 = ~n7959 & n7962;
  assign n7964 = n7959 & ~n7962;
  assign n7965 = ~n7963 & ~n7964;
  assign n7966 = ~n7946 & ~n7953;
  assign n7967 = ~n7965 & n7966;
  assign n7968 = ~n7959 & ~n7962;
  assign n7969 = ~n7967 & ~n7968;
  assign n7970 = ~n7963 & n7966;
  assign n7971 = ~n7964 & n7970;
  assign n7972 = ~n7965 & ~n7966;
  assign n7973 = ~n7971 & ~n7972;
  assign n7974 = ~n7969 & ~n7973;
  assign n7975 = ~n7956 & ~n7974;
  assign n7976 = ~A79  & A80 ;
  assign n7977 = A79  & ~A80 ;
  assign n7978 = A81  & ~n7977;
  assign n7979 = ~n7976 & n7978;
  assign n7980 = ~n7976 & ~n7977;
  assign n7981 = ~A81  & ~n7980;
  assign n7982 = ~n7979 & ~n7981;
  assign n7983 = ~A82  & A83 ;
  assign n7984 = A82  & ~A83 ;
  assign n7985 = A84  & ~n7984;
  assign n7986 = ~n7983 & n7985;
  assign n7987 = ~n7983 & ~n7984;
  assign n7988 = ~A84  & ~n7987;
  assign n7989 = ~n7986 & ~n7988;
  assign n7990 = ~n7982 & n7989;
  assign n7991 = n7982 & ~n7989;
  assign n7992 = ~n7990 & ~n7991;
  assign n7993 = A82  & A83 ;
  assign n7994 = A84  & ~n7987;
  assign n7995 = ~n7993 & ~n7994;
  assign n7996 = A79  & A80 ;
  assign n7997 = A81  & ~n7980;
  assign n7998 = ~n7996 & ~n7997;
  assign n7999 = ~n7995 & n7998;
  assign n8000 = n7995 & ~n7998;
  assign n8001 = ~n7999 & ~n8000;
  assign n8002 = ~n7982 & ~n7989;
  assign n8003 = ~n8001 & n8002;
  assign n8004 = ~n7995 & ~n7998;
  assign n8005 = ~n8003 & ~n8004;
  assign n8006 = ~n7999 & n8002;
  assign n8007 = ~n8000 & n8006;
  assign n8008 = ~n8001 & ~n8002;
  assign n8009 = ~n8007 & ~n8008;
  assign n8010 = ~n8005 & ~n8009;
  assign n8011 = ~n7992 & ~n8010;
  assign n8012 = ~n7975 & n8011;
  assign n8013 = n7975 & ~n8011;
  assign n8014 = ~n8012 & ~n8013;
  assign n8015 = ~n7939 & n8014;
  assign n8016 = n7939 & ~n8014;
  assign n8017 = ~n8015 & ~n8016;
  assign n8018 = ~n7864 & n8017;
  assign n8019 = n7864 & ~n8017;
  assign n8020 = ~n8018 & ~n8019;
  assign n8021 = ~n7711 & n8020;
  assign n8022 = n7711 & ~n8020;
  assign n8023 = ~n8021 & ~n8022;
  assign n8024 = ~n7402 & ~n8023;
  assign n8025 = ~n7399 & n8024;
  assign n8026 = ~n7394 & n8025;
  assign n8027 = ~n7394 & ~n7399;
  assign n8028 = ~n8024 & ~n8027;
  assign n8029 = ~n8026 & ~n8028;
  assign n8030 = ~n7608 & ~n7621;
  assign n8031 = ~n7625 & ~n8030;
  assign n8032 = ~n7572 & ~n7608;
  assign n8033 = ~n7590 & n8032;
  assign n8034 = ~n7626 & n8033;
  assign n8035 = ~n7572 & ~n7585;
  assign n8036 = ~n7589 & ~n8035;
  assign n8037 = ~n8034 & ~n8036;
  assign n8038 = ~n7589 & n8032;
  assign n8039 = ~n7590 & n8038;
  assign n8040 = ~n7626 & ~n8035;
  assign n8041 = n8039 & n8040;
  assign n8042 = ~n8037 & ~n8041;
  assign n8043 = n8031 & ~n8042;
  assign n8044 = ~n8034 & n8036;
  assign n8045 = n8034 & ~n8036;
  assign n8046 = ~n8044 & ~n8045;
  assign n8047 = ~n8031 & ~n8046;
  assign n8048 = ~n7630 & ~n7705;
  assign n8049 = ~n8047 & n8048;
  assign n8050 = ~n8043 & n8049;
  assign n8051 = ~n8043 & ~n8047;
  assign n8052 = ~n8048 & ~n8051;
  assign n8053 = ~n8050 & ~n8052;
  assign n8054 = ~n7683 & ~n7696;
  assign n8055 = ~n7700 & ~n8054;
  assign n8056 = ~n7647 & ~n7683;
  assign n8057 = ~n7665 & n8056;
  assign n8058 = ~n7701 & n8057;
  assign n8059 = ~n7647 & ~n7660;
  assign n8060 = ~n7664 & ~n8059;
  assign n8061 = ~n8058 & n8060;
  assign n8062 = n8058 & ~n8060;
  assign n8063 = ~n8061 & ~n8062;
  assign n8064 = ~n8055 & ~n8063;
  assign n8065 = ~n8058 & ~n8060;
  assign n8066 = ~n7664 & n8056;
  assign n8067 = ~n7665 & n8066;
  assign n8068 = ~n7701 & ~n8059;
  assign n8069 = n8067 & n8068;
  assign n8070 = ~n8065 & ~n8069;
  assign n8071 = n8055 & ~n8070;
  assign n8072 = ~n8064 & ~n8071;
  assign n8073 = ~n8053 & n8072;
  assign n8074 = ~n8047 & ~n8048;
  assign n8075 = ~n8043 & n8074;
  assign n8076 = n8048 & ~n8051;
  assign n8077 = ~n8075 & ~n8076;
  assign n8078 = ~n8072 & ~n8077;
  assign n8079 = ~n8073 & ~n8078;
  assign n8080 = ~n7530 & ~n7543;
  assign n8081 = ~n7547 & ~n8080;
  assign n8082 = ~n7494 & ~n7530;
  assign n8083 = ~n7512 & n8082;
  assign n8084 = ~n7548 & n8083;
  assign n8085 = ~n7494 & ~n7507;
  assign n8086 = ~n7511 & ~n8085;
  assign n8087 = ~n8084 & n8086;
  assign n8088 = n8084 & ~n8086;
  assign n8089 = ~n8087 & ~n8088;
  assign n8090 = ~n8081 & ~n8089;
  assign n8091 = ~n8084 & ~n8086;
  assign n8092 = ~n7511 & n8082;
  assign n8093 = ~n7512 & n8092;
  assign n8094 = ~n7548 & ~n8085;
  assign n8095 = n8093 & n8094;
  assign n8096 = ~n8091 & ~n8095;
  assign n8097 = n8081 & ~n8096;
  assign n8098 = ~n8090 & ~n8097;
  assign n8099 = ~n7455 & ~n7468;
  assign n8100 = ~n7472 & ~n8099;
  assign n8101 = ~n7419 & ~n7455;
  assign n8102 = ~n7437 & n8101;
  assign n8103 = ~n7473 & n8102;
  assign n8104 = ~n7419 & ~n7432;
  assign n8105 = ~n7436 & ~n8104;
  assign n8106 = ~n8103 & ~n8105;
  assign n8107 = ~n7436 & n8101;
  assign n8108 = ~n7437 & n8107;
  assign n8109 = ~n7473 & ~n8104;
  assign n8110 = n8108 & n8109;
  assign n8111 = ~n8106 & ~n8110;
  assign n8112 = n8100 & ~n8111;
  assign n8113 = ~n8103 & n8105;
  assign n8114 = n8103 & ~n8105;
  assign n8115 = ~n8113 & ~n8114;
  assign n8116 = ~n8100 & ~n8115;
  assign n8117 = ~n7477 & ~n7552;
  assign n8118 = ~n8116 & ~n8117;
  assign n8119 = ~n8112 & n8118;
  assign n8120 = ~n8112 & ~n8116;
  assign n8121 = n8117 & ~n8120;
  assign n8122 = ~n8119 & ~n8121;
  assign n8123 = ~n8098 & ~n8122;
  assign n8124 = ~n8116 & n8117;
  assign n8125 = ~n8112 & n8124;
  assign n8126 = ~n8117 & ~n8120;
  assign n8127 = ~n8125 & ~n8126;
  assign n8128 = n8098 & ~n8127;
  assign n8129 = ~n7555 & ~n7708;
  assign n8130 = ~n8128 & ~n8129;
  assign n8131 = ~n8123 & n8130;
  assign n8132 = ~n8123 & ~n8128;
  assign n8133 = n8129 & ~n8132;
  assign n8134 = ~n8131 & ~n8133;
  assign n8135 = ~n8079 & ~n8134;
  assign n8136 = ~n8128 & n8129;
  assign n8137 = ~n8123 & n8136;
  assign n8138 = ~n8129 & ~n8132;
  assign n8139 = ~n8137 & ~n8138;
  assign n8140 = n8079 & ~n8139;
  assign n8141 = ~n7711 & ~n8020;
  assign n8142 = ~n8140 & n8141;
  assign n8143 = ~n8135 & n8142;
  assign n8144 = ~n8135 & ~n8140;
  assign n8145 = ~n8141 & ~n8144;
  assign n8146 = ~n8143 & ~n8145;
  assign n8147 = ~n7839 & ~n7852;
  assign n8148 = ~n7856 & ~n8147;
  assign n8149 = ~n7803 & ~n7839;
  assign n8150 = ~n7821 & n8149;
  assign n8151 = ~n7857 & n8150;
  assign n8152 = ~n7803 & ~n7816;
  assign n8153 = ~n7820 & ~n8152;
  assign n8154 = ~n8151 & n8153;
  assign n8155 = n8151 & ~n8153;
  assign n8156 = ~n8154 & ~n8155;
  assign n8157 = ~n8148 & ~n8156;
  assign n8158 = ~n8151 & ~n8153;
  assign n8159 = ~n7820 & n8149;
  assign n8160 = ~n7821 & n8159;
  assign n8161 = ~n7857 & ~n8152;
  assign n8162 = n8160 & n8161;
  assign n8163 = ~n8158 & ~n8162;
  assign n8164 = n8148 & ~n8163;
  assign n8165 = ~n8157 & ~n8164;
  assign n8166 = ~n7764 & ~n7777;
  assign n8167 = ~n7781 & ~n8166;
  assign n8168 = ~n7728 & ~n7764;
  assign n8169 = ~n7746 & n8168;
  assign n8170 = ~n7782 & n8169;
  assign n8171 = ~n7728 & ~n7741;
  assign n8172 = ~n7745 & ~n8171;
  assign n8173 = ~n8170 & ~n8172;
  assign n8174 = ~n7745 & n8168;
  assign n8175 = ~n7746 & n8174;
  assign n8176 = ~n7782 & ~n8171;
  assign n8177 = n8175 & n8176;
  assign n8178 = ~n8173 & ~n8177;
  assign n8179 = n8167 & ~n8178;
  assign n8180 = ~n8170 & n8172;
  assign n8181 = n8170 & ~n8172;
  assign n8182 = ~n8180 & ~n8181;
  assign n8183 = ~n8167 & ~n8182;
  assign n8184 = ~n7786 & ~n7861;
  assign n8185 = ~n8183 & ~n8184;
  assign n8186 = ~n8179 & n8185;
  assign n8187 = ~n8179 & ~n8183;
  assign n8188 = n8184 & ~n8187;
  assign n8189 = ~n8186 & ~n8188;
  assign n8190 = ~n8165 & ~n8189;
  assign n8191 = ~n8183 & n8184;
  assign n8192 = ~n8179 & n8191;
  assign n8193 = ~n8184 & ~n8187;
  assign n8194 = ~n8192 & ~n8193;
  assign n8195 = n8165 & ~n8194;
  assign n8196 = ~n7864 & ~n8017;
  assign n8197 = ~n8195 & n8196;
  assign n8198 = ~n8190 & n8197;
  assign n8199 = ~n8190 & ~n8195;
  assign n8200 = ~n8196 & ~n8199;
  assign n8201 = ~n8198 & ~n8200;
  assign n8202 = ~n7917 & ~n7930;
  assign n8203 = ~n7934 & ~n8202;
  assign n8204 = ~n7881 & ~n7917;
  assign n8205 = ~n7899 & n8204;
  assign n8206 = ~n7935 & n8205;
  assign n8207 = ~n7881 & ~n7894;
  assign n8208 = ~n7898 & ~n8207;
  assign n8209 = ~n8206 & ~n8208;
  assign n8210 = ~n7898 & n8204;
  assign n8211 = ~n7899 & n8210;
  assign n8212 = ~n7935 & ~n8207;
  assign n8213 = n8211 & n8212;
  assign n8214 = ~n8209 & ~n8213;
  assign n8215 = n8203 & ~n8214;
  assign n8216 = ~n8206 & n8208;
  assign n8217 = n8206 & ~n8208;
  assign n8218 = ~n8216 & ~n8217;
  assign n8219 = ~n8203 & ~n8218;
  assign n8220 = ~n7939 & ~n8014;
  assign n8221 = ~n8219 & n8220;
  assign n8222 = ~n8215 & n8221;
  assign n8223 = ~n8215 & ~n8219;
  assign n8224 = ~n8220 & ~n8223;
  assign n8225 = ~n8222 & ~n8224;
  assign n8226 = ~n7992 & ~n8005;
  assign n8227 = ~n8009 & ~n8226;
  assign n8228 = ~n7956 & ~n7992;
  assign n8229 = ~n7974 & n8228;
  assign n8230 = ~n8010 & n8229;
  assign n8231 = ~n7956 & ~n7969;
  assign n8232 = ~n7973 & ~n8231;
  assign n8233 = ~n8230 & n8232;
  assign n8234 = n8230 & ~n8232;
  assign n8235 = ~n8233 & ~n8234;
  assign n8236 = ~n8227 & ~n8235;
  assign n8237 = ~n8230 & ~n8232;
  assign n8238 = ~n7973 & n8228;
  assign n8239 = ~n7974 & n8238;
  assign n8240 = ~n8010 & ~n8231;
  assign n8241 = n8239 & n8240;
  assign n8242 = ~n8237 & ~n8241;
  assign n8243 = n8227 & ~n8242;
  assign n8244 = ~n8236 & ~n8243;
  assign n8245 = ~n8225 & n8244;
  assign n8246 = ~n8219 & ~n8220;
  assign n8247 = ~n8215 & n8246;
  assign n8248 = n8220 & ~n8223;
  assign n8249 = ~n8247 & ~n8248;
  assign n8250 = ~n8244 & ~n8249;
  assign n8251 = ~n8245 & ~n8250;
  assign n8252 = ~n8201 & n8251;
  assign n8253 = ~n8195 & ~n8196;
  assign n8254 = ~n8190 & n8253;
  assign n8255 = n8196 & ~n8199;
  assign n8256 = ~n8254 & ~n8255;
  assign n8257 = ~n8251 & ~n8256;
  assign n8258 = ~n8252 & ~n8257;
  assign n8259 = ~n8146 & n8258;
  assign n8260 = ~n8140 & ~n8141;
  assign n8261 = ~n8135 & n8260;
  assign n8262 = n8141 & ~n8144;
  assign n8263 = ~n8261 & ~n8262;
  assign n8264 = ~n8258 & ~n8263;
  assign n8265 = ~n8259 & ~n8264;
  assign n8266 = ~n8029 & n8265;
  assign n8267 = ~n7399 & ~n8024;
  assign n8268 = ~n7394 & n8267;
  assign n8269 = n8024 & ~n8027;
  assign n8270 = ~n8268 & ~n8269;
  assign n8271 = ~n8265 & ~n8270;
  assign n8272 = ~n8266 & ~n8271;
  assign n8273 = A334  & A335 ;
  assign n8274 = A334  & ~A335 ;
  assign n8275 = ~A334  & A335 ;
  assign n8276 = ~n8274 & ~n8275;
  assign n8277 = A336  & ~n8276;
  assign n8278 = ~n8273 & ~n8277;
  assign n8279 = A331  & A332 ;
  assign n8280 = A331  & ~A332 ;
  assign n8281 = ~A331  & A332 ;
  assign n8282 = ~n8280 & ~n8281;
  assign n8283 = A333  & ~n8282;
  assign n8284 = ~n8279 & ~n8283;
  assign n8285 = n8278 & ~n8284;
  assign n8286 = ~n8278 & n8284;
  assign n8287 = A333  & ~n8280;
  assign n8288 = ~n8281 & n8287;
  assign n8289 = ~A333  & ~n8282;
  assign n8290 = ~n8288 & ~n8289;
  assign n8291 = A336  & ~n8274;
  assign n8292 = ~n8275 & n8291;
  assign n8293 = ~A336  & ~n8276;
  assign n8294 = ~n8292 & ~n8293;
  assign n8295 = ~n8290 & ~n8294;
  assign n8296 = ~n8286 & n8295;
  assign n8297 = ~n8285 & n8296;
  assign n8298 = ~n8285 & ~n8286;
  assign n8299 = ~n8295 & ~n8298;
  assign n8300 = ~n8297 & ~n8299;
  assign n8301 = ~n8290 & n8294;
  assign n8302 = n8290 & ~n8294;
  assign n8303 = ~n8301 & ~n8302;
  assign n8304 = n8295 & ~n8298;
  assign n8305 = ~n8278 & ~n8284;
  assign n8306 = ~n8304 & ~n8305;
  assign n8307 = ~n8303 & ~n8306;
  assign n8308 = ~n8300 & ~n8307;
  assign n8309 = ~n8300 & ~n8306;
  assign n8310 = A340  & A341 ;
  assign n8311 = A340  & ~A341 ;
  assign n8312 = ~A340  & A341 ;
  assign n8313 = ~n8311 & ~n8312;
  assign n8314 = A342  & ~n8313;
  assign n8315 = ~n8310 & ~n8314;
  assign n8316 = A337  & A338 ;
  assign n8317 = A337  & ~A338 ;
  assign n8318 = ~A337  & A338 ;
  assign n8319 = ~n8317 & ~n8318;
  assign n8320 = A339  & ~n8319;
  assign n8321 = ~n8316 & ~n8320;
  assign n8322 = ~n8315 & n8321;
  assign n8323 = n8315 & ~n8321;
  assign n8324 = ~n8322 & ~n8323;
  assign n8325 = A339  & ~n8317;
  assign n8326 = ~n8318 & n8325;
  assign n8327 = ~A339  & ~n8319;
  assign n8328 = ~n8326 & ~n8327;
  assign n8329 = A342  & ~n8311;
  assign n8330 = ~n8312 & n8329;
  assign n8331 = ~A342  & ~n8313;
  assign n8332 = ~n8330 & ~n8331;
  assign n8333 = ~n8328 & ~n8332;
  assign n8334 = ~n8324 & n8333;
  assign n8335 = ~n8315 & ~n8321;
  assign n8336 = ~n8334 & ~n8335;
  assign n8337 = ~n8322 & n8333;
  assign n8338 = ~n8323 & n8337;
  assign n8339 = ~n8324 & ~n8333;
  assign n8340 = ~n8338 & ~n8339;
  assign n8341 = ~n8336 & ~n8340;
  assign n8342 = ~n8328 & n8332;
  assign n8343 = n8328 & ~n8332;
  assign n8344 = ~n8342 & ~n8343;
  assign n8345 = ~n8303 & ~n8344;
  assign n8346 = ~n8341 & n8345;
  assign n8347 = ~n8309 & n8346;
  assign n8348 = ~n8336 & ~n8344;
  assign n8349 = ~n8340 & ~n8348;
  assign n8350 = ~n8347 & ~n8349;
  assign n8351 = ~n8340 & n8345;
  assign n8352 = ~n8341 & n8351;
  assign n8353 = ~n8309 & ~n8348;
  assign n8354 = n8352 & n8353;
  assign n8355 = ~n8350 & ~n8354;
  assign n8356 = n8308 & ~n8355;
  assign n8357 = ~n8347 & n8349;
  assign n8358 = n8347 & ~n8349;
  assign n8359 = ~n8357 & ~n8358;
  assign n8360 = ~n8308 & ~n8359;
  assign n8361 = ~n8341 & ~n8344;
  assign n8362 = ~n8303 & ~n8309;
  assign n8363 = ~n8361 & n8362;
  assign n8364 = n8361 & ~n8362;
  assign n8365 = ~n8363 & ~n8364;
  assign n8366 = ~A325  & A326 ;
  assign n8367 = A325  & ~A326 ;
  assign n8368 = A327  & ~n8367;
  assign n8369 = ~n8366 & n8368;
  assign n8370 = ~n8366 & ~n8367;
  assign n8371 = ~A327  & ~n8370;
  assign n8372 = ~n8369 & ~n8371;
  assign n8373 = ~A328  & A329 ;
  assign n8374 = A328  & ~A329 ;
  assign n8375 = A330  & ~n8374;
  assign n8376 = ~n8373 & n8375;
  assign n8377 = ~n8373 & ~n8374;
  assign n8378 = ~A330  & ~n8377;
  assign n8379 = ~n8376 & ~n8378;
  assign n8380 = ~n8372 & n8379;
  assign n8381 = n8372 & ~n8379;
  assign n8382 = ~n8380 & ~n8381;
  assign n8383 = A328  & A329 ;
  assign n8384 = A330  & ~n8377;
  assign n8385 = ~n8383 & ~n8384;
  assign n8386 = A325  & A326 ;
  assign n8387 = A327  & ~n8370;
  assign n8388 = ~n8386 & ~n8387;
  assign n8389 = ~n8385 & n8388;
  assign n8390 = n8385 & ~n8388;
  assign n8391 = ~n8389 & ~n8390;
  assign n8392 = ~n8372 & ~n8379;
  assign n8393 = ~n8391 & n8392;
  assign n8394 = ~n8385 & ~n8388;
  assign n8395 = ~n8393 & ~n8394;
  assign n8396 = ~n8389 & n8392;
  assign n8397 = ~n8390 & n8396;
  assign n8398 = ~n8391 & ~n8392;
  assign n8399 = ~n8397 & ~n8398;
  assign n8400 = ~n8395 & ~n8399;
  assign n8401 = ~n8382 & ~n8400;
  assign n8402 = ~A319  & A320 ;
  assign n8403 = A319  & ~A320 ;
  assign n8404 = A321  & ~n8403;
  assign n8405 = ~n8402 & n8404;
  assign n8406 = ~n8402 & ~n8403;
  assign n8407 = ~A321  & ~n8406;
  assign n8408 = ~n8405 & ~n8407;
  assign n8409 = ~A322  & A323 ;
  assign n8410 = A322  & ~A323 ;
  assign n8411 = A324  & ~n8410;
  assign n8412 = ~n8409 & n8411;
  assign n8413 = ~n8409 & ~n8410;
  assign n8414 = ~A324  & ~n8413;
  assign n8415 = ~n8412 & ~n8414;
  assign n8416 = ~n8408 & n8415;
  assign n8417 = n8408 & ~n8415;
  assign n8418 = ~n8416 & ~n8417;
  assign n8419 = A322  & A323 ;
  assign n8420 = A324  & ~n8413;
  assign n8421 = ~n8419 & ~n8420;
  assign n8422 = A319  & A320 ;
  assign n8423 = A321  & ~n8406;
  assign n8424 = ~n8422 & ~n8423;
  assign n8425 = ~n8421 & n8424;
  assign n8426 = n8421 & ~n8424;
  assign n8427 = ~n8425 & ~n8426;
  assign n8428 = ~n8408 & ~n8415;
  assign n8429 = ~n8427 & n8428;
  assign n8430 = ~n8421 & ~n8424;
  assign n8431 = ~n8429 & ~n8430;
  assign n8432 = ~n8425 & n8428;
  assign n8433 = ~n8426 & n8432;
  assign n8434 = ~n8427 & ~n8428;
  assign n8435 = ~n8433 & ~n8434;
  assign n8436 = ~n8431 & ~n8435;
  assign n8437 = ~n8418 & ~n8436;
  assign n8438 = ~n8401 & n8437;
  assign n8439 = n8401 & ~n8437;
  assign n8440 = ~n8438 & ~n8439;
  assign n8441 = ~n8365 & ~n8440;
  assign n8442 = ~n8360 & n8441;
  assign n8443 = ~n8356 & n8442;
  assign n8444 = ~n8356 & ~n8360;
  assign n8445 = ~n8441 & ~n8444;
  assign n8446 = ~n8443 & ~n8445;
  assign n8447 = ~n8418 & ~n8431;
  assign n8448 = ~n8435 & ~n8447;
  assign n8449 = ~n8382 & ~n8418;
  assign n8450 = ~n8400 & n8449;
  assign n8451 = ~n8436 & n8450;
  assign n8452 = ~n8382 & ~n8395;
  assign n8453 = ~n8399 & ~n8452;
  assign n8454 = ~n8451 & n8453;
  assign n8455 = n8451 & ~n8453;
  assign n8456 = ~n8454 & ~n8455;
  assign n8457 = ~n8448 & ~n8456;
  assign n8458 = ~n8451 & ~n8453;
  assign n8459 = ~n8399 & n8449;
  assign n8460 = ~n8400 & n8459;
  assign n8461 = ~n8436 & ~n8452;
  assign n8462 = n8460 & n8461;
  assign n8463 = ~n8458 & ~n8462;
  assign n8464 = n8448 & ~n8463;
  assign n8465 = ~n8457 & ~n8464;
  assign n8466 = ~n8446 & n8465;
  assign n8467 = ~n8360 & ~n8441;
  assign n8468 = ~n8356 & n8467;
  assign n8469 = n8441 & ~n8444;
  assign n8470 = ~n8468 & ~n8469;
  assign n8471 = ~n8465 & ~n8470;
  assign n8472 = ~n8466 & ~n8471;
  assign n8473 = A346  & A347 ;
  assign n8474 = A346  & ~A347 ;
  assign n8475 = ~A346  & A347 ;
  assign n8476 = ~n8474 & ~n8475;
  assign n8477 = A348  & ~n8476;
  assign n8478 = ~n8473 & ~n8477;
  assign n8479 = A343  & A344 ;
  assign n8480 = A343  & ~A344 ;
  assign n8481 = ~A343  & A344 ;
  assign n8482 = ~n8480 & ~n8481;
  assign n8483 = A345  & ~n8482;
  assign n8484 = ~n8479 & ~n8483;
  assign n8485 = n8478 & ~n8484;
  assign n8486 = ~n8478 & n8484;
  assign n8487 = A345  & ~n8480;
  assign n8488 = ~n8481 & n8487;
  assign n8489 = ~A345  & ~n8482;
  assign n8490 = ~n8488 & ~n8489;
  assign n8491 = A348  & ~n8474;
  assign n8492 = ~n8475 & n8491;
  assign n8493 = ~A348  & ~n8476;
  assign n8494 = ~n8492 & ~n8493;
  assign n8495 = ~n8490 & ~n8494;
  assign n8496 = ~n8486 & n8495;
  assign n8497 = ~n8485 & n8496;
  assign n8498 = ~n8485 & ~n8486;
  assign n8499 = ~n8495 & ~n8498;
  assign n8500 = ~n8497 & ~n8499;
  assign n8501 = ~n8490 & n8494;
  assign n8502 = n8490 & ~n8494;
  assign n8503 = ~n8501 & ~n8502;
  assign n8504 = n8495 & ~n8498;
  assign n8505 = ~n8478 & ~n8484;
  assign n8506 = ~n8504 & ~n8505;
  assign n8507 = ~n8503 & ~n8506;
  assign n8508 = ~n8500 & ~n8507;
  assign n8509 = ~n8500 & ~n8506;
  assign n8510 = A352  & A353 ;
  assign n8511 = A352  & ~A353 ;
  assign n8512 = ~A352  & A353 ;
  assign n8513 = ~n8511 & ~n8512;
  assign n8514 = A354  & ~n8513;
  assign n8515 = ~n8510 & ~n8514;
  assign n8516 = A349  & A350 ;
  assign n8517 = A349  & ~A350 ;
  assign n8518 = ~A349  & A350 ;
  assign n8519 = ~n8517 & ~n8518;
  assign n8520 = A351  & ~n8519;
  assign n8521 = ~n8516 & ~n8520;
  assign n8522 = ~n8515 & n8521;
  assign n8523 = n8515 & ~n8521;
  assign n8524 = ~n8522 & ~n8523;
  assign n8525 = A351  & ~n8517;
  assign n8526 = ~n8518 & n8525;
  assign n8527 = ~A351  & ~n8519;
  assign n8528 = ~n8526 & ~n8527;
  assign n8529 = A354  & ~n8511;
  assign n8530 = ~n8512 & n8529;
  assign n8531 = ~A354  & ~n8513;
  assign n8532 = ~n8530 & ~n8531;
  assign n8533 = ~n8528 & ~n8532;
  assign n8534 = ~n8524 & n8533;
  assign n8535 = ~n8515 & ~n8521;
  assign n8536 = ~n8534 & ~n8535;
  assign n8537 = ~n8522 & n8533;
  assign n8538 = ~n8523 & n8537;
  assign n8539 = ~n8524 & ~n8533;
  assign n8540 = ~n8538 & ~n8539;
  assign n8541 = ~n8536 & ~n8540;
  assign n8542 = ~n8528 & n8532;
  assign n8543 = n8528 & ~n8532;
  assign n8544 = ~n8542 & ~n8543;
  assign n8545 = ~n8503 & ~n8544;
  assign n8546 = ~n8541 & n8545;
  assign n8547 = ~n8509 & n8546;
  assign n8548 = ~n8536 & ~n8544;
  assign n8549 = ~n8540 & ~n8548;
  assign n8550 = ~n8547 & n8549;
  assign n8551 = n8547 & ~n8549;
  assign n8552 = ~n8550 & ~n8551;
  assign n8553 = ~n8508 & ~n8552;
  assign n8554 = ~n8547 & ~n8549;
  assign n8555 = ~n8540 & n8545;
  assign n8556 = ~n8541 & n8555;
  assign n8557 = ~n8509 & ~n8548;
  assign n8558 = n8556 & n8557;
  assign n8559 = ~n8554 & ~n8558;
  assign n8560 = n8508 & ~n8559;
  assign n8561 = ~n8553 & ~n8560;
  assign n8562 = A358  & A359 ;
  assign n8563 = A358  & ~A359 ;
  assign n8564 = ~A358  & A359 ;
  assign n8565 = ~n8563 & ~n8564;
  assign n8566 = A360  & ~n8565;
  assign n8567 = ~n8562 & ~n8566;
  assign n8568 = A355  & A356 ;
  assign n8569 = A355  & ~A356 ;
  assign n8570 = ~A355  & A356 ;
  assign n8571 = ~n8569 & ~n8570;
  assign n8572 = A357  & ~n8571;
  assign n8573 = ~n8568 & ~n8572;
  assign n8574 = n8567 & ~n8573;
  assign n8575 = ~n8567 & n8573;
  assign n8576 = A357  & ~n8569;
  assign n8577 = ~n8570 & n8576;
  assign n8578 = ~A357  & ~n8571;
  assign n8579 = ~n8577 & ~n8578;
  assign n8580 = A360  & ~n8563;
  assign n8581 = ~n8564 & n8580;
  assign n8582 = ~A360  & ~n8565;
  assign n8583 = ~n8581 & ~n8582;
  assign n8584 = ~n8579 & ~n8583;
  assign n8585 = ~n8575 & n8584;
  assign n8586 = ~n8574 & n8585;
  assign n8587 = ~n8574 & ~n8575;
  assign n8588 = ~n8584 & ~n8587;
  assign n8589 = ~n8586 & ~n8588;
  assign n8590 = ~n8579 & n8583;
  assign n8591 = n8579 & ~n8583;
  assign n8592 = ~n8590 & ~n8591;
  assign n8593 = n8584 & ~n8587;
  assign n8594 = ~n8567 & ~n8573;
  assign n8595 = ~n8593 & ~n8594;
  assign n8596 = ~n8592 & ~n8595;
  assign n8597 = ~n8589 & ~n8596;
  assign n8598 = ~n8589 & ~n8595;
  assign n8599 = A364  & A365 ;
  assign n8600 = A364  & ~A365 ;
  assign n8601 = ~A364  & A365 ;
  assign n8602 = ~n8600 & ~n8601;
  assign n8603 = A366  & ~n8602;
  assign n8604 = ~n8599 & ~n8603;
  assign n8605 = A361  & A362 ;
  assign n8606 = A361  & ~A362 ;
  assign n8607 = ~A361  & A362 ;
  assign n8608 = ~n8606 & ~n8607;
  assign n8609 = A363  & ~n8608;
  assign n8610 = ~n8605 & ~n8609;
  assign n8611 = ~n8604 & n8610;
  assign n8612 = n8604 & ~n8610;
  assign n8613 = ~n8611 & ~n8612;
  assign n8614 = A363  & ~n8606;
  assign n8615 = ~n8607 & n8614;
  assign n8616 = ~A363  & ~n8608;
  assign n8617 = ~n8615 & ~n8616;
  assign n8618 = A366  & ~n8600;
  assign n8619 = ~n8601 & n8618;
  assign n8620 = ~A366  & ~n8602;
  assign n8621 = ~n8619 & ~n8620;
  assign n8622 = ~n8617 & ~n8621;
  assign n8623 = ~n8613 & n8622;
  assign n8624 = ~n8604 & ~n8610;
  assign n8625 = ~n8623 & ~n8624;
  assign n8626 = ~n8611 & n8622;
  assign n8627 = ~n8612 & n8626;
  assign n8628 = ~n8613 & ~n8622;
  assign n8629 = ~n8627 & ~n8628;
  assign n8630 = ~n8625 & ~n8629;
  assign n8631 = ~n8617 & n8621;
  assign n8632 = n8617 & ~n8621;
  assign n8633 = ~n8631 & ~n8632;
  assign n8634 = ~n8592 & ~n8633;
  assign n8635 = ~n8630 & n8634;
  assign n8636 = ~n8598 & n8635;
  assign n8637 = ~n8625 & ~n8633;
  assign n8638 = ~n8629 & ~n8637;
  assign n8639 = ~n8636 & ~n8638;
  assign n8640 = ~n8629 & n8634;
  assign n8641 = ~n8630 & n8640;
  assign n8642 = ~n8598 & ~n8637;
  assign n8643 = n8641 & n8642;
  assign n8644 = ~n8639 & ~n8643;
  assign n8645 = n8597 & ~n8644;
  assign n8646 = ~n8636 & n8638;
  assign n8647 = n8636 & ~n8638;
  assign n8648 = ~n8646 & ~n8647;
  assign n8649 = ~n8597 & ~n8648;
  assign n8650 = ~n8630 & ~n8633;
  assign n8651 = ~n8592 & ~n8598;
  assign n8652 = ~n8650 & n8651;
  assign n8653 = n8650 & ~n8651;
  assign n8654 = ~n8652 & ~n8653;
  assign n8655 = ~n8541 & ~n8544;
  assign n8656 = ~n8503 & ~n8509;
  assign n8657 = ~n8655 & n8656;
  assign n8658 = n8655 & ~n8656;
  assign n8659 = ~n8657 & ~n8658;
  assign n8660 = ~n8654 & ~n8659;
  assign n8661 = ~n8649 & ~n8660;
  assign n8662 = ~n8645 & n8661;
  assign n8663 = ~n8645 & ~n8649;
  assign n8664 = n8660 & ~n8663;
  assign n8665 = ~n8662 & ~n8664;
  assign n8666 = ~n8561 & ~n8665;
  assign n8667 = ~n8649 & n8660;
  assign n8668 = ~n8645 & n8667;
  assign n8669 = ~n8660 & ~n8663;
  assign n8670 = ~n8668 & ~n8669;
  assign n8671 = n8561 & ~n8670;
  assign n8672 = ~n8654 & n8659;
  assign n8673 = n8654 & ~n8659;
  assign n8674 = ~n8672 & ~n8673;
  assign n8675 = ~n8365 & n8440;
  assign n8676 = n8365 & ~n8440;
  assign n8677 = ~n8675 & ~n8676;
  assign n8678 = ~n8674 & ~n8677;
  assign n8679 = ~n8671 & ~n8678;
  assign n8680 = ~n8666 & n8679;
  assign n8681 = ~n8666 & ~n8671;
  assign n8682 = n8678 & ~n8681;
  assign n8683 = ~n8680 & ~n8682;
  assign n8684 = ~n8472 & ~n8683;
  assign n8685 = ~n8671 & n8678;
  assign n8686 = ~n8666 & n8685;
  assign n8687 = ~n8678 & ~n8681;
  assign n8688 = ~n8686 & ~n8687;
  assign n8689 = n8472 & ~n8688;
  assign n8690 = ~n8674 & n8677;
  assign n8691 = n8674 & ~n8677;
  assign n8692 = ~n8690 & ~n8691;
  assign n8693 = ~A313  & A314 ;
  assign n8694 = A313  & ~A314 ;
  assign n8695 = A315  & ~n8694;
  assign n8696 = ~n8693 & n8695;
  assign n8697 = ~n8693 & ~n8694;
  assign n8698 = ~A315  & ~n8697;
  assign n8699 = ~n8696 & ~n8698;
  assign n8700 = ~A316  & A317 ;
  assign n8701 = A316  & ~A317 ;
  assign n8702 = A318  & ~n8701;
  assign n8703 = ~n8700 & n8702;
  assign n8704 = ~n8700 & ~n8701;
  assign n8705 = ~A318  & ~n8704;
  assign n8706 = ~n8703 & ~n8705;
  assign n8707 = ~n8699 & n8706;
  assign n8708 = n8699 & ~n8706;
  assign n8709 = ~n8707 & ~n8708;
  assign n8710 = A316  & A317 ;
  assign n8711 = A318  & ~n8704;
  assign n8712 = ~n8710 & ~n8711;
  assign n8713 = A313  & A314 ;
  assign n8714 = A315  & ~n8697;
  assign n8715 = ~n8713 & ~n8714;
  assign n8716 = ~n8712 & n8715;
  assign n8717 = n8712 & ~n8715;
  assign n8718 = ~n8716 & ~n8717;
  assign n8719 = ~n8699 & ~n8706;
  assign n8720 = ~n8718 & n8719;
  assign n8721 = ~n8712 & ~n8715;
  assign n8722 = ~n8720 & ~n8721;
  assign n8723 = ~n8716 & n8719;
  assign n8724 = ~n8717 & n8723;
  assign n8725 = ~n8718 & ~n8719;
  assign n8726 = ~n8724 & ~n8725;
  assign n8727 = ~n8722 & ~n8726;
  assign n8728 = ~n8709 & ~n8727;
  assign n8729 = ~A307  & A308 ;
  assign n8730 = A307  & ~A308 ;
  assign n8731 = A309  & ~n8730;
  assign n8732 = ~n8729 & n8731;
  assign n8733 = ~n8729 & ~n8730;
  assign n8734 = ~A309  & ~n8733;
  assign n8735 = ~n8732 & ~n8734;
  assign n8736 = ~A310  & A311 ;
  assign n8737 = A310  & ~A311 ;
  assign n8738 = A312  & ~n8737;
  assign n8739 = ~n8736 & n8738;
  assign n8740 = ~n8736 & ~n8737;
  assign n8741 = ~A312  & ~n8740;
  assign n8742 = ~n8739 & ~n8741;
  assign n8743 = ~n8735 & n8742;
  assign n8744 = n8735 & ~n8742;
  assign n8745 = ~n8743 & ~n8744;
  assign n8746 = A310  & A311 ;
  assign n8747 = A312  & ~n8740;
  assign n8748 = ~n8746 & ~n8747;
  assign n8749 = A307  & A308 ;
  assign n8750 = A309  & ~n8733;
  assign n8751 = ~n8749 & ~n8750;
  assign n8752 = ~n8748 & n8751;
  assign n8753 = n8748 & ~n8751;
  assign n8754 = ~n8752 & ~n8753;
  assign n8755 = ~n8735 & ~n8742;
  assign n8756 = ~n8754 & n8755;
  assign n8757 = ~n8748 & ~n8751;
  assign n8758 = ~n8756 & ~n8757;
  assign n8759 = ~n8752 & n8755;
  assign n8760 = ~n8753 & n8759;
  assign n8761 = ~n8754 & ~n8755;
  assign n8762 = ~n8760 & ~n8761;
  assign n8763 = ~n8758 & ~n8762;
  assign n8764 = ~n8745 & ~n8763;
  assign n8765 = ~n8728 & n8764;
  assign n8766 = n8728 & ~n8764;
  assign n8767 = ~n8765 & ~n8766;
  assign n8768 = ~A301  & A302 ;
  assign n8769 = A301  & ~A302 ;
  assign n8770 = A303  & ~n8769;
  assign n8771 = ~n8768 & n8770;
  assign n8772 = ~n8768 & ~n8769;
  assign n8773 = ~A303  & ~n8772;
  assign n8774 = ~n8771 & ~n8773;
  assign n8775 = ~A304  & A305 ;
  assign n8776 = A304  & ~A305 ;
  assign n8777 = A306  & ~n8776;
  assign n8778 = ~n8775 & n8777;
  assign n8779 = ~n8775 & ~n8776;
  assign n8780 = ~A306  & ~n8779;
  assign n8781 = ~n8778 & ~n8780;
  assign n8782 = ~n8774 & n8781;
  assign n8783 = n8774 & ~n8781;
  assign n8784 = ~n8782 & ~n8783;
  assign n8785 = A304  & A305 ;
  assign n8786 = A306  & ~n8779;
  assign n8787 = ~n8785 & ~n8786;
  assign n8788 = A301  & A302 ;
  assign n8789 = A303  & ~n8772;
  assign n8790 = ~n8788 & ~n8789;
  assign n8791 = ~n8787 & n8790;
  assign n8792 = n8787 & ~n8790;
  assign n8793 = ~n8791 & ~n8792;
  assign n8794 = ~n8774 & ~n8781;
  assign n8795 = ~n8793 & n8794;
  assign n8796 = ~n8787 & ~n8790;
  assign n8797 = ~n8795 & ~n8796;
  assign n8798 = ~n8791 & n8794;
  assign n8799 = ~n8792 & n8798;
  assign n8800 = ~n8793 & ~n8794;
  assign n8801 = ~n8799 & ~n8800;
  assign n8802 = ~n8797 & ~n8801;
  assign n8803 = ~n8784 & ~n8802;
  assign n8804 = ~A295  & A296 ;
  assign n8805 = A295  & ~A296 ;
  assign n8806 = A297  & ~n8805;
  assign n8807 = ~n8804 & n8806;
  assign n8808 = ~n8804 & ~n8805;
  assign n8809 = ~A297  & ~n8808;
  assign n8810 = ~n8807 & ~n8809;
  assign n8811 = ~A298  & A299 ;
  assign n8812 = A298  & ~A299 ;
  assign n8813 = A300  & ~n8812;
  assign n8814 = ~n8811 & n8813;
  assign n8815 = ~n8811 & ~n8812;
  assign n8816 = ~A300  & ~n8815;
  assign n8817 = ~n8814 & ~n8816;
  assign n8818 = ~n8810 & n8817;
  assign n8819 = n8810 & ~n8817;
  assign n8820 = ~n8818 & ~n8819;
  assign n8821 = A298  & A299 ;
  assign n8822 = A300  & ~n8815;
  assign n8823 = ~n8821 & ~n8822;
  assign n8824 = A295  & A296 ;
  assign n8825 = A297  & ~n8808;
  assign n8826 = ~n8824 & ~n8825;
  assign n8827 = ~n8823 & n8826;
  assign n8828 = n8823 & ~n8826;
  assign n8829 = ~n8827 & ~n8828;
  assign n8830 = ~n8810 & ~n8817;
  assign n8831 = ~n8829 & n8830;
  assign n8832 = ~n8823 & ~n8826;
  assign n8833 = ~n8831 & ~n8832;
  assign n8834 = ~n8827 & n8830;
  assign n8835 = ~n8828 & n8834;
  assign n8836 = ~n8829 & ~n8830;
  assign n8837 = ~n8835 & ~n8836;
  assign n8838 = ~n8833 & ~n8837;
  assign n8839 = ~n8820 & ~n8838;
  assign n8840 = ~n8803 & n8839;
  assign n8841 = n8803 & ~n8839;
  assign n8842 = ~n8840 & ~n8841;
  assign n8843 = ~n8767 & n8842;
  assign n8844 = n8767 & ~n8842;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = ~A289  & A290 ;
  assign n8847 = A289  & ~A290 ;
  assign n8848 = A291  & ~n8847;
  assign n8849 = ~n8846 & n8848;
  assign n8850 = ~n8846 & ~n8847;
  assign n8851 = ~A291  & ~n8850;
  assign n8852 = ~n8849 & ~n8851;
  assign n8853 = ~A292  & A293 ;
  assign n8854 = A292  & ~A293 ;
  assign n8855 = A294  & ~n8854;
  assign n8856 = ~n8853 & n8855;
  assign n8857 = ~n8853 & ~n8854;
  assign n8858 = ~A294  & ~n8857;
  assign n8859 = ~n8856 & ~n8858;
  assign n8860 = ~n8852 & n8859;
  assign n8861 = n8852 & ~n8859;
  assign n8862 = ~n8860 & ~n8861;
  assign n8863 = A292  & A293 ;
  assign n8864 = A294  & ~n8857;
  assign n8865 = ~n8863 & ~n8864;
  assign n8866 = A289  & A290 ;
  assign n8867 = A291  & ~n8850;
  assign n8868 = ~n8866 & ~n8867;
  assign n8869 = ~n8865 & n8868;
  assign n8870 = n8865 & ~n8868;
  assign n8871 = ~n8869 & ~n8870;
  assign n8872 = ~n8852 & ~n8859;
  assign n8873 = ~n8871 & n8872;
  assign n8874 = ~n8865 & ~n8868;
  assign n8875 = ~n8873 & ~n8874;
  assign n8876 = ~n8869 & n8872;
  assign n8877 = ~n8870 & n8876;
  assign n8878 = ~n8871 & ~n8872;
  assign n8879 = ~n8877 & ~n8878;
  assign n8880 = ~n8875 & ~n8879;
  assign n8881 = ~n8862 & ~n8880;
  assign n8882 = ~A283  & A284 ;
  assign n8883 = A283  & ~A284 ;
  assign n8884 = A285  & ~n8883;
  assign n8885 = ~n8882 & n8884;
  assign n8886 = ~n8882 & ~n8883;
  assign n8887 = ~A285  & ~n8886;
  assign n8888 = ~n8885 & ~n8887;
  assign n8889 = ~A286  & A287 ;
  assign n8890 = A286  & ~A287 ;
  assign n8891 = A288  & ~n8890;
  assign n8892 = ~n8889 & n8891;
  assign n8893 = ~n8889 & ~n8890;
  assign n8894 = ~A288  & ~n8893;
  assign n8895 = ~n8892 & ~n8894;
  assign n8896 = ~n8888 & n8895;
  assign n8897 = n8888 & ~n8895;
  assign n8898 = ~n8896 & ~n8897;
  assign n8899 = A286  & A287 ;
  assign n8900 = A288  & ~n8893;
  assign n8901 = ~n8899 & ~n8900;
  assign n8902 = A283  & A284 ;
  assign n8903 = A285  & ~n8886;
  assign n8904 = ~n8902 & ~n8903;
  assign n8905 = ~n8901 & n8904;
  assign n8906 = n8901 & ~n8904;
  assign n8907 = ~n8905 & ~n8906;
  assign n8908 = ~n8888 & ~n8895;
  assign n8909 = ~n8907 & n8908;
  assign n8910 = ~n8901 & ~n8904;
  assign n8911 = ~n8909 & ~n8910;
  assign n8912 = ~n8905 & n8908;
  assign n8913 = ~n8906 & n8912;
  assign n8914 = ~n8907 & ~n8908;
  assign n8915 = ~n8913 & ~n8914;
  assign n8916 = ~n8911 & ~n8915;
  assign n8917 = ~n8898 & ~n8916;
  assign n8918 = ~n8881 & n8917;
  assign n8919 = n8881 & ~n8917;
  assign n8920 = ~n8918 & ~n8919;
  assign n8921 = ~A277  & A278 ;
  assign n8922 = A277  & ~A278 ;
  assign n8923 = A279  & ~n8922;
  assign n8924 = ~n8921 & n8923;
  assign n8925 = ~n8921 & ~n8922;
  assign n8926 = ~A279  & ~n8925;
  assign n8927 = ~n8924 & ~n8926;
  assign n8928 = ~A280  & A281 ;
  assign n8929 = A280  & ~A281 ;
  assign n8930 = A282  & ~n8929;
  assign n8931 = ~n8928 & n8930;
  assign n8932 = ~n8928 & ~n8929;
  assign n8933 = ~A282  & ~n8932;
  assign n8934 = ~n8931 & ~n8933;
  assign n8935 = ~n8927 & n8934;
  assign n8936 = n8927 & ~n8934;
  assign n8937 = ~n8935 & ~n8936;
  assign n8938 = A280  & A281 ;
  assign n8939 = A282  & ~n8932;
  assign n8940 = ~n8938 & ~n8939;
  assign n8941 = A277  & A278 ;
  assign n8942 = A279  & ~n8925;
  assign n8943 = ~n8941 & ~n8942;
  assign n8944 = ~n8940 & n8943;
  assign n8945 = n8940 & ~n8943;
  assign n8946 = ~n8944 & ~n8945;
  assign n8947 = ~n8927 & ~n8934;
  assign n8948 = ~n8946 & n8947;
  assign n8949 = ~n8940 & ~n8943;
  assign n8950 = ~n8948 & ~n8949;
  assign n8951 = ~n8944 & n8947;
  assign n8952 = ~n8945 & n8951;
  assign n8953 = ~n8946 & ~n8947;
  assign n8954 = ~n8952 & ~n8953;
  assign n8955 = ~n8950 & ~n8954;
  assign n8956 = ~n8937 & ~n8955;
  assign n8957 = ~A271  & A272 ;
  assign n8958 = A271  & ~A272 ;
  assign n8959 = A273  & ~n8958;
  assign n8960 = ~n8957 & n8959;
  assign n8961 = ~n8957 & ~n8958;
  assign n8962 = ~A273  & ~n8961;
  assign n8963 = ~n8960 & ~n8962;
  assign n8964 = ~A274  & A275 ;
  assign n8965 = A274  & ~A275 ;
  assign n8966 = A276  & ~n8965;
  assign n8967 = ~n8964 & n8966;
  assign n8968 = ~n8964 & ~n8965;
  assign n8969 = ~A276  & ~n8968;
  assign n8970 = ~n8967 & ~n8969;
  assign n8971 = ~n8963 & n8970;
  assign n8972 = n8963 & ~n8970;
  assign n8973 = ~n8971 & ~n8972;
  assign n8974 = A274  & A275 ;
  assign n8975 = A276  & ~n8968;
  assign n8976 = ~n8974 & ~n8975;
  assign n8977 = A271  & A272 ;
  assign n8978 = A273  & ~n8961;
  assign n8979 = ~n8977 & ~n8978;
  assign n8980 = ~n8976 & n8979;
  assign n8981 = n8976 & ~n8979;
  assign n8982 = ~n8980 & ~n8981;
  assign n8983 = ~n8963 & ~n8970;
  assign n8984 = ~n8982 & n8983;
  assign n8985 = ~n8976 & ~n8979;
  assign n8986 = ~n8984 & ~n8985;
  assign n8987 = ~n8980 & n8983;
  assign n8988 = ~n8981 & n8987;
  assign n8989 = ~n8982 & ~n8983;
  assign n8990 = ~n8988 & ~n8989;
  assign n8991 = ~n8986 & ~n8990;
  assign n8992 = ~n8973 & ~n8991;
  assign n8993 = ~n8956 & n8992;
  assign n8994 = n8956 & ~n8992;
  assign n8995 = ~n8993 & ~n8994;
  assign n8996 = ~n8920 & n8995;
  assign n8997 = n8920 & ~n8995;
  assign n8998 = ~n8996 & ~n8997;
  assign n8999 = ~n8845 & n8998;
  assign n9000 = n8845 & ~n8998;
  assign n9001 = ~n8999 & ~n9000;
  assign n9002 = ~n8692 & ~n9001;
  assign n9003 = ~n8689 & n9002;
  assign n9004 = ~n8684 & n9003;
  assign n9005 = ~n8684 & ~n8689;
  assign n9006 = ~n9002 & ~n9005;
  assign n9007 = ~n9004 & ~n9006;
  assign n9008 = ~n8820 & ~n8833;
  assign n9009 = ~n8837 & ~n9008;
  assign n9010 = ~n8784 & ~n8820;
  assign n9011 = ~n8802 & n9010;
  assign n9012 = ~n8838 & n9011;
  assign n9013 = ~n8784 & ~n8797;
  assign n9014 = ~n8801 & ~n9013;
  assign n9015 = ~n9012 & n9014;
  assign n9016 = n9012 & ~n9014;
  assign n9017 = ~n9015 & ~n9016;
  assign n9018 = ~n9009 & ~n9017;
  assign n9019 = ~n9012 & ~n9014;
  assign n9020 = ~n8801 & n9010;
  assign n9021 = ~n8802 & n9020;
  assign n9022 = ~n8838 & ~n9013;
  assign n9023 = n9021 & n9022;
  assign n9024 = ~n9019 & ~n9023;
  assign n9025 = n9009 & ~n9024;
  assign n9026 = ~n9018 & ~n9025;
  assign n9027 = ~n8745 & ~n8758;
  assign n9028 = ~n8762 & ~n9027;
  assign n9029 = ~n8709 & ~n8745;
  assign n9030 = ~n8727 & n9029;
  assign n9031 = ~n8763 & n9030;
  assign n9032 = ~n8709 & ~n8722;
  assign n9033 = ~n8726 & ~n9032;
  assign n9034 = ~n9031 & ~n9033;
  assign n9035 = ~n8726 & n9029;
  assign n9036 = ~n8727 & n9035;
  assign n9037 = ~n8763 & ~n9032;
  assign n9038 = n9036 & n9037;
  assign n9039 = ~n9034 & ~n9038;
  assign n9040 = n9028 & ~n9039;
  assign n9041 = ~n9031 & n9033;
  assign n9042 = n9031 & ~n9033;
  assign n9043 = ~n9041 & ~n9042;
  assign n9044 = ~n9028 & ~n9043;
  assign n9045 = ~n8767 & ~n8842;
  assign n9046 = ~n9044 & ~n9045;
  assign n9047 = ~n9040 & n9046;
  assign n9048 = ~n9040 & ~n9044;
  assign n9049 = n9045 & ~n9048;
  assign n9050 = ~n9047 & ~n9049;
  assign n9051 = ~n9026 & ~n9050;
  assign n9052 = ~n9044 & n9045;
  assign n9053 = ~n9040 & n9052;
  assign n9054 = ~n9045 & ~n9048;
  assign n9055 = ~n9053 & ~n9054;
  assign n9056 = n9026 & ~n9055;
  assign n9057 = ~n8845 & ~n8998;
  assign n9058 = ~n9056 & n9057;
  assign n9059 = ~n9051 & n9058;
  assign n9060 = ~n9051 & ~n9056;
  assign n9061 = ~n9057 & ~n9060;
  assign n9062 = ~n9059 & ~n9061;
  assign n9063 = ~n8898 & ~n8911;
  assign n9064 = ~n8915 & ~n9063;
  assign n9065 = ~n8862 & ~n8898;
  assign n9066 = ~n8880 & n9065;
  assign n9067 = ~n8916 & n9066;
  assign n9068 = ~n8862 & ~n8875;
  assign n9069 = ~n8879 & ~n9068;
  assign n9070 = ~n9067 & ~n9069;
  assign n9071 = ~n8879 & n9065;
  assign n9072 = ~n8880 & n9071;
  assign n9073 = ~n8916 & ~n9068;
  assign n9074 = n9072 & n9073;
  assign n9075 = ~n9070 & ~n9074;
  assign n9076 = n9064 & ~n9075;
  assign n9077 = ~n9067 & n9069;
  assign n9078 = n9067 & ~n9069;
  assign n9079 = ~n9077 & ~n9078;
  assign n9080 = ~n9064 & ~n9079;
  assign n9081 = ~n8920 & ~n8995;
  assign n9082 = ~n9080 & n9081;
  assign n9083 = ~n9076 & n9082;
  assign n9084 = ~n9076 & ~n9080;
  assign n9085 = ~n9081 & ~n9084;
  assign n9086 = ~n9083 & ~n9085;
  assign n9087 = ~n8973 & ~n8986;
  assign n9088 = ~n8990 & ~n9087;
  assign n9089 = ~n8937 & ~n8973;
  assign n9090 = ~n8955 & n9089;
  assign n9091 = ~n8991 & n9090;
  assign n9092 = ~n8937 & ~n8950;
  assign n9093 = ~n8954 & ~n9092;
  assign n9094 = ~n9091 & n9093;
  assign n9095 = n9091 & ~n9093;
  assign n9096 = ~n9094 & ~n9095;
  assign n9097 = ~n9088 & ~n9096;
  assign n9098 = ~n9091 & ~n9093;
  assign n9099 = ~n8954 & n9089;
  assign n9100 = ~n8955 & n9099;
  assign n9101 = ~n8991 & ~n9092;
  assign n9102 = n9100 & n9101;
  assign n9103 = ~n9098 & ~n9102;
  assign n9104 = n9088 & ~n9103;
  assign n9105 = ~n9097 & ~n9104;
  assign n9106 = ~n9086 & n9105;
  assign n9107 = ~n9080 & ~n9081;
  assign n9108 = ~n9076 & n9107;
  assign n9109 = n9081 & ~n9084;
  assign n9110 = ~n9108 & ~n9109;
  assign n9111 = ~n9105 & ~n9110;
  assign n9112 = ~n9106 & ~n9111;
  assign n9113 = ~n9062 & n9112;
  assign n9114 = ~n9056 & ~n9057;
  assign n9115 = ~n9051 & n9114;
  assign n9116 = n9057 & ~n9060;
  assign n9117 = ~n9115 & ~n9116;
  assign n9118 = ~n9112 & ~n9117;
  assign n9119 = ~n9113 & ~n9118;
  assign n9120 = ~n9007 & n9119;
  assign n9121 = ~n8689 & ~n9002;
  assign n9122 = ~n8684 & n9121;
  assign n9123 = n9002 & ~n9005;
  assign n9124 = ~n9122 & ~n9123;
  assign n9125 = ~n9119 & ~n9124;
  assign n9126 = ~n9120 & ~n9125;
  assign n9127 = A394  & A395 ;
  assign n9128 = A394  & ~A395 ;
  assign n9129 = ~A394  & A395 ;
  assign n9130 = ~n9128 & ~n9129;
  assign n9131 = A396  & ~n9130;
  assign n9132 = ~n9127 & ~n9131;
  assign n9133 = A391  & A392 ;
  assign n9134 = A391  & ~A392 ;
  assign n9135 = ~A391  & A392 ;
  assign n9136 = ~n9134 & ~n9135;
  assign n9137 = A393  & ~n9136;
  assign n9138 = ~n9133 & ~n9137;
  assign n9139 = n9132 & ~n9138;
  assign n9140 = ~n9132 & n9138;
  assign n9141 = A393  & ~n9134;
  assign n9142 = ~n9135 & n9141;
  assign n9143 = ~A393  & ~n9136;
  assign n9144 = ~n9142 & ~n9143;
  assign n9145 = A396  & ~n9128;
  assign n9146 = ~n9129 & n9145;
  assign n9147 = ~A396  & ~n9130;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = ~n9144 & ~n9148;
  assign n9150 = ~n9140 & n9149;
  assign n9151 = ~n9139 & n9150;
  assign n9152 = ~n9139 & ~n9140;
  assign n9153 = ~n9149 & ~n9152;
  assign n9154 = ~n9151 & ~n9153;
  assign n9155 = ~n9144 & n9148;
  assign n9156 = n9144 & ~n9148;
  assign n9157 = ~n9155 & ~n9156;
  assign n9158 = n9149 & ~n9152;
  assign n9159 = ~n9132 & ~n9138;
  assign n9160 = ~n9158 & ~n9159;
  assign n9161 = ~n9157 & ~n9160;
  assign n9162 = ~n9154 & ~n9161;
  assign n9163 = ~n9154 & ~n9160;
  assign n9164 = A400  & A401 ;
  assign n9165 = A400  & ~A401 ;
  assign n9166 = ~A400  & A401 ;
  assign n9167 = ~n9165 & ~n9166;
  assign n9168 = A402  & ~n9167;
  assign n9169 = ~n9164 & ~n9168;
  assign n9170 = A397  & A398 ;
  assign n9171 = A397  & ~A398 ;
  assign n9172 = ~A397  & A398 ;
  assign n9173 = ~n9171 & ~n9172;
  assign n9174 = A399  & ~n9173;
  assign n9175 = ~n9170 & ~n9174;
  assign n9176 = ~n9169 & n9175;
  assign n9177 = n9169 & ~n9175;
  assign n9178 = ~n9176 & ~n9177;
  assign n9179 = A399  & ~n9171;
  assign n9180 = ~n9172 & n9179;
  assign n9181 = ~A399  & ~n9173;
  assign n9182 = ~n9180 & ~n9181;
  assign n9183 = A402  & ~n9165;
  assign n9184 = ~n9166 & n9183;
  assign n9185 = ~A402  & ~n9167;
  assign n9186 = ~n9184 & ~n9185;
  assign n9187 = ~n9182 & ~n9186;
  assign n9188 = ~n9178 & n9187;
  assign n9189 = ~n9169 & ~n9175;
  assign n9190 = ~n9188 & ~n9189;
  assign n9191 = ~n9176 & n9187;
  assign n9192 = ~n9177 & n9191;
  assign n9193 = ~n9178 & ~n9187;
  assign n9194 = ~n9192 & ~n9193;
  assign n9195 = ~n9190 & ~n9194;
  assign n9196 = ~n9182 & n9186;
  assign n9197 = n9182 & ~n9186;
  assign n9198 = ~n9196 & ~n9197;
  assign n9199 = ~n9157 & ~n9198;
  assign n9200 = ~n9195 & n9199;
  assign n9201 = ~n9163 & n9200;
  assign n9202 = ~n9190 & ~n9198;
  assign n9203 = ~n9194 & ~n9202;
  assign n9204 = ~n9201 & n9203;
  assign n9205 = n9201 & ~n9203;
  assign n9206 = ~n9204 & ~n9205;
  assign n9207 = ~n9162 & ~n9206;
  assign n9208 = ~n9201 & ~n9203;
  assign n9209 = ~n9194 & n9199;
  assign n9210 = ~n9195 & n9209;
  assign n9211 = ~n9163 & ~n9202;
  assign n9212 = n9210 & n9211;
  assign n9213 = ~n9208 & ~n9212;
  assign n9214 = n9162 & ~n9213;
  assign n9215 = ~n9207 & ~n9214;
  assign n9216 = A406  & A407 ;
  assign n9217 = A406  & ~A407 ;
  assign n9218 = ~A406  & A407 ;
  assign n9219 = ~n9217 & ~n9218;
  assign n9220 = A408  & ~n9219;
  assign n9221 = ~n9216 & ~n9220;
  assign n9222 = A403  & A404 ;
  assign n9223 = A403  & ~A404 ;
  assign n9224 = ~A403  & A404 ;
  assign n9225 = ~n9223 & ~n9224;
  assign n9226 = A405  & ~n9225;
  assign n9227 = ~n9222 & ~n9226;
  assign n9228 = n9221 & ~n9227;
  assign n9229 = ~n9221 & n9227;
  assign n9230 = A405  & ~n9223;
  assign n9231 = ~n9224 & n9230;
  assign n9232 = ~A405  & ~n9225;
  assign n9233 = ~n9231 & ~n9232;
  assign n9234 = A408  & ~n9217;
  assign n9235 = ~n9218 & n9234;
  assign n9236 = ~A408  & ~n9219;
  assign n9237 = ~n9235 & ~n9236;
  assign n9238 = ~n9233 & ~n9237;
  assign n9239 = ~n9229 & n9238;
  assign n9240 = ~n9228 & n9239;
  assign n9241 = ~n9228 & ~n9229;
  assign n9242 = ~n9238 & ~n9241;
  assign n9243 = ~n9240 & ~n9242;
  assign n9244 = ~n9233 & n9237;
  assign n9245 = n9233 & ~n9237;
  assign n9246 = ~n9244 & ~n9245;
  assign n9247 = n9238 & ~n9241;
  assign n9248 = ~n9221 & ~n9227;
  assign n9249 = ~n9247 & ~n9248;
  assign n9250 = ~n9246 & ~n9249;
  assign n9251 = ~n9243 & ~n9250;
  assign n9252 = ~n9243 & ~n9249;
  assign n9253 = A412  & A413 ;
  assign n9254 = A412  & ~A413 ;
  assign n9255 = ~A412  & A413 ;
  assign n9256 = ~n9254 & ~n9255;
  assign n9257 = A414  & ~n9256;
  assign n9258 = ~n9253 & ~n9257;
  assign n9259 = A409  & A410 ;
  assign n9260 = A409  & ~A410 ;
  assign n9261 = ~A409  & A410 ;
  assign n9262 = ~n9260 & ~n9261;
  assign n9263 = A411  & ~n9262;
  assign n9264 = ~n9259 & ~n9263;
  assign n9265 = ~n9258 & n9264;
  assign n9266 = n9258 & ~n9264;
  assign n9267 = ~n9265 & ~n9266;
  assign n9268 = A411  & ~n9260;
  assign n9269 = ~n9261 & n9268;
  assign n9270 = ~A411  & ~n9262;
  assign n9271 = ~n9269 & ~n9270;
  assign n9272 = A414  & ~n9254;
  assign n9273 = ~n9255 & n9272;
  assign n9274 = ~A414  & ~n9256;
  assign n9275 = ~n9273 & ~n9274;
  assign n9276 = ~n9271 & ~n9275;
  assign n9277 = ~n9267 & n9276;
  assign n9278 = ~n9258 & ~n9264;
  assign n9279 = ~n9277 & ~n9278;
  assign n9280 = ~n9265 & n9276;
  assign n9281 = ~n9266 & n9280;
  assign n9282 = ~n9267 & ~n9276;
  assign n9283 = ~n9281 & ~n9282;
  assign n9284 = ~n9279 & ~n9283;
  assign n9285 = ~n9271 & n9275;
  assign n9286 = n9271 & ~n9275;
  assign n9287 = ~n9285 & ~n9286;
  assign n9288 = ~n9246 & ~n9287;
  assign n9289 = ~n9284 & n9288;
  assign n9290 = ~n9252 & n9289;
  assign n9291 = ~n9279 & ~n9287;
  assign n9292 = ~n9283 & ~n9291;
  assign n9293 = ~n9290 & ~n9292;
  assign n9294 = ~n9283 & n9288;
  assign n9295 = ~n9284 & n9294;
  assign n9296 = ~n9252 & ~n9291;
  assign n9297 = n9295 & n9296;
  assign n9298 = ~n9293 & ~n9297;
  assign n9299 = n9251 & ~n9298;
  assign n9300 = ~n9290 & n9292;
  assign n9301 = n9290 & ~n9292;
  assign n9302 = ~n9300 & ~n9301;
  assign n9303 = ~n9251 & ~n9302;
  assign n9304 = ~n9284 & ~n9287;
  assign n9305 = ~n9246 & ~n9252;
  assign n9306 = ~n9304 & n9305;
  assign n9307 = n9304 & ~n9305;
  assign n9308 = ~n9306 & ~n9307;
  assign n9309 = ~n9195 & ~n9198;
  assign n9310 = ~n9157 & ~n9163;
  assign n9311 = ~n9309 & n9310;
  assign n9312 = n9309 & ~n9310;
  assign n9313 = ~n9311 & ~n9312;
  assign n9314 = ~n9308 & ~n9313;
  assign n9315 = ~n9303 & ~n9314;
  assign n9316 = ~n9299 & n9315;
  assign n9317 = ~n9299 & ~n9303;
  assign n9318 = n9314 & ~n9317;
  assign n9319 = ~n9316 & ~n9318;
  assign n9320 = ~n9215 & ~n9319;
  assign n9321 = ~n9303 & n9314;
  assign n9322 = ~n9299 & n9321;
  assign n9323 = ~n9314 & ~n9317;
  assign n9324 = ~n9322 & ~n9323;
  assign n9325 = n9215 & ~n9324;
  assign n9326 = ~n9308 & n9313;
  assign n9327 = n9308 & ~n9313;
  assign n9328 = ~n9326 & ~n9327;
  assign n9329 = ~A385  & A386 ;
  assign n9330 = A385  & ~A386 ;
  assign n9331 = A387  & ~n9330;
  assign n9332 = ~n9329 & n9331;
  assign n9333 = ~n9329 & ~n9330;
  assign n9334 = ~A387  & ~n9333;
  assign n9335 = ~n9332 & ~n9334;
  assign n9336 = ~A388  & A389 ;
  assign n9337 = A388  & ~A389 ;
  assign n9338 = A390  & ~n9337;
  assign n9339 = ~n9336 & n9338;
  assign n9340 = ~n9336 & ~n9337;
  assign n9341 = ~A390  & ~n9340;
  assign n9342 = ~n9339 & ~n9341;
  assign n9343 = ~n9335 & n9342;
  assign n9344 = n9335 & ~n9342;
  assign n9345 = ~n9343 & ~n9344;
  assign n9346 = A388  & A389 ;
  assign n9347 = A390  & ~n9340;
  assign n9348 = ~n9346 & ~n9347;
  assign n9349 = A385  & A386 ;
  assign n9350 = A387  & ~n9333;
  assign n9351 = ~n9349 & ~n9350;
  assign n9352 = ~n9348 & n9351;
  assign n9353 = n9348 & ~n9351;
  assign n9354 = ~n9352 & ~n9353;
  assign n9355 = ~n9335 & ~n9342;
  assign n9356 = ~n9354 & n9355;
  assign n9357 = ~n9348 & ~n9351;
  assign n9358 = ~n9356 & ~n9357;
  assign n9359 = ~n9352 & n9355;
  assign n9360 = ~n9353 & n9359;
  assign n9361 = ~n9354 & ~n9355;
  assign n9362 = ~n9360 & ~n9361;
  assign n9363 = ~n9358 & ~n9362;
  assign n9364 = ~n9345 & ~n9363;
  assign n9365 = ~A379  & A380 ;
  assign n9366 = A379  & ~A380 ;
  assign n9367 = A381  & ~n9366;
  assign n9368 = ~n9365 & n9367;
  assign n9369 = ~n9365 & ~n9366;
  assign n9370 = ~A381  & ~n9369;
  assign n9371 = ~n9368 & ~n9370;
  assign n9372 = ~A382  & A383 ;
  assign n9373 = A382  & ~A383 ;
  assign n9374 = A384  & ~n9373;
  assign n9375 = ~n9372 & n9374;
  assign n9376 = ~n9372 & ~n9373;
  assign n9377 = ~A384  & ~n9376;
  assign n9378 = ~n9375 & ~n9377;
  assign n9379 = ~n9371 & n9378;
  assign n9380 = n9371 & ~n9378;
  assign n9381 = ~n9379 & ~n9380;
  assign n9382 = A382  & A383 ;
  assign n9383 = A384  & ~n9376;
  assign n9384 = ~n9382 & ~n9383;
  assign n9385 = A379  & A380 ;
  assign n9386 = A381  & ~n9369;
  assign n9387 = ~n9385 & ~n9386;
  assign n9388 = ~n9384 & n9387;
  assign n9389 = n9384 & ~n9387;
  assign n9390 = ~n9388 & ~n9389;
  assign n9391 = ~n9371 & ~n9378;
  assign n9392 = ~n9390 & n9391;
  assign n9393 = ~n9384 & ~n9387;
  assign n9394 = ~n9392 & ~n9393;
  assign n9395 = ~n9388 & n9391;
  assign n9396 = ~n9389 & n9395;
  assign n9397 = ~n9390 & ~n9391;
  assign n9398 = ~n9396 & ~n9397;
  assign n9399 = ~n9394 & ~n9398;
  assign n9400 = ~n9381 & ~n9399;
  assign n9401 = ~n9364 & n9400;
  assign n9402 = n9364 & ~n9400;
  assign n9403 = ~n9401 & ~n9402;
  assign n9404 = ~A373  & A374 ;
  assign n9405 = A373  & ~A374 ;
  assign n9406 = A375  & ~n9405;
  assign n9407 = ~n9404 & n9406;
  assign n9408 = ~n9404 & ~n9405;
  assign n9409 = ~A375  & ~n9408;
  assign n9410 = ~n9407 & ~n9409;
  assign n9411 = ~A376  & A377 ;
  assign n9412 = A376  & ~A377 ;
  assign n9413 = A378  & ~n9412;
  assign n9414 = ~n9411 & n9413;
  assign n9415 = ~n9411 & ~n9412;
  assign n9416 = ~A378  & ~n9415;
  assign n9417 = ~n9414 & ~n9416;
  assign n9418 = ~n9410 & n9417;
  assign n9419 = n9410 & ~n9417;
  assign n9420 = ~n9418 & ~n9419;
  assign n9421 = A376  & A377 ;
  assign n9422 = A378  & ~n9415;
  assign n9423 = ~n9421 & ~n9422;
  assign n9424 = A373  & A374 ;
  assign n9425 = A375  & ~n9408;
  assign n9426 = ~n9424 & ~n9425;
  assign n9427 = ~n9423 & n9426;
  assign n9428 = n9423 & ~n9426;
  assign n9429 = ~n9427 & ~n9428;
  assign n9430 = ~n9410 & ~n9417;
  assign n9431 = ~n9429 & n9430;
  assign n9432 = ~n9423 & ~n9426;
  assign n9433 = ~n9431 & ~n9432;
  assign n9434 = ~n9427 & n9430;
  assign n9435 = ~n9428 & n9434;
  assign n9436 = ~n9429 & ~n9430;
  assign n9437 = ~n9435 & ~n9436;
  assign n9438 = ~n9433 & ~n9437;
  assign n9439 = ~n9420 & ~n9438;
  assign n9440 = ~A367  & A368 ;
  assign n9441 = A367  & ~A368 ;
  assign n9442 = A369  & ~n9441;
  assign n9443 = ~n9440 & n9442;
  assign n9444 = ~n9440 & ~n9441;
  assign n9445 = ~A369  & ~n9444;
  assign n9446 = ~n9443 & ~n9445;
  assign n9447 = ~A370  & A371 ;
  assign n9448 = A370  & ~A371 ;
  assign n9449 = A372  & ~n9448;
  assign n9450 = ~n9447 & n9449;
  assign n9451 = ~n9447 & ~n9448;
  assign n9452 = ~A372  & ~n9451;
  assign n9453 = ~n9450 & ~n9452;
  assign n9454 = ~n9446 & n9453;
  assign n9455 = n9446 & ~n9453;
  assign n9456 = ~n9454 & ~n9455;
  assign n9457 = A370  & A371 ;
  assign n9458 = A372  & ~n9451;
  assign n9459 = ~n9457 & ~n9458;
  assign n9460 = A367  & A368 ;
  assign n9461 = A369  & ~n9444;
  assign n9462 = ~n9460 & ~n9461;
  assign n9463 = ~n9459 & n9462;
  assign n9464 = n9459 & ~n9462;
  assign n9465 = ~n9463 & ~n9464;
  assign n9466 = ~n9446 & ~n9453;
  assign n9467 = ~n9465 & n9466;
  assign n9468 = ~n9459 & ~n9462;
  assign n9469 = ~n9467 & ~n9468;
  assign n9470 = ~n9463 & n9466;
  assign n9471 = ~n9464 & n9470;
  assign n9472 = ~n9465 & ~n9466;
  assign n9473 = ~n9471 & ~n9472;
  assign n9474 = ~n9469 & ~n9473;
  assign n9475 = ~n9456 & ~n9474;
  assign n9476 = ~n9439 & n9475;
  assign n9477 = n9439 & ~n9475;
  assign n9478 = ~n9476 & ~n9477;
  assign n9479 = ~n9403 & n9478;
  assign n9480 = n9403 & ~n9478;
  assign n9481 = ~n9479 & ~n9480;
  assign n9482 = ~n9328 & ~n9481;
  assign n9483 = ~n9325 & n9482;
  assign n9484 = ~n9320 & n9483;
  assign n9485 = ~n9320 & ~n9325;
  assign n9486 = ~n9482 & ~n9485;
  assign n9487 = ~n9484 & ~n9486;
  assign n9488 = ~n9381 & ~n9394;
  assign n9489 = ~n9398 & ~n9488;
  assign n9490 = ~n9345 & ~n9381;
  assign n9491 = ~n9363 & n9490;
  assign n9492 = ~n9399 & n9491;
  assign n9493 = ~n9345 & ~n9358;
  assign n9494 = ~n9362 & ~n9493;
  assign n9495 = ~n9492 & ~n9494;
  assign n9496 = ~n9362 & n9490;
  assign n9497 = ~n9363 & n9496;
  assign n9498 = ~n9399 & ~n9493;
  assign n9499 = n9497 & n9498;
  assign n9500 = ~n9495 & ~n9499;
  assign n9501 = n9489 & ~n9500;
  assign n9502 = ~n9492 & n9494;
  assign n9503 = n9492 & ~n9494;
  assign n9504 = ~n9502 & ~n9503;
  assign n9505 = ~n9489 & ~n9504;
  assign n9506 = ~n9403 & ~n9478;
  assign n9507 = ~n9505 & n9506;
  assign n9508 = ~n9501 & n9507;
  assign n9509 = ~n9501 & ~n9505;
  assign n9510 = ~n9506 & ~n9509;
  assign n9511 = ~n9508 & ~n9510;
  assign n9512 = ~n9456 & ~n9469;
  assign n9513 = ~n9473 & ~n9512;
  assign n9514 = ~n9420 & ~n9456;
  assign n9515 = ~n9438 & n9514;
  assign n9516 = ~n9474 & n9515;
  assign n9517 = ~n9420 & ~n9433;
  assign n9518 = ~n9437 & ~n9517;
  assign n9519 = ~n9516 & n9518;
  assign n9520 = n9516 & ~n9518;
  assign n9521 = ~n9519 & ~n9520;
  assign n9522 = ~n9513 & ~n9521;
  assign n9523 = ~n9516 & ~n9518;
  assign n9524 = ~n9437 & n9514;
  assign n9525 = ~n9438 & n9524;
  assign n9526 = ~n9474 & ~n9517;
  assign n9527 = n9525 & n9526;
  assign n9528 = ~n9523 & ~n9527;
  assign n9529 = n9513 & ~n9528;
  assign n9530 = ~n9522 & ~n9529;
  assign n9531 = ~n9511 & n9530;
  assign n9532 = ~n9505 & ~n9506;
  assign n9533 = ~n9501 & n9532;
  assign n9534 = n9506 & ~n9509;
  assign n9535 = ~n9533 & ~n9534;
  assign n9536 = ~n9530 & ~n9535;
  assign n9537 = ~n9531 & ~n9536;
  assign n9538 = ~n9487 & n9537;
  assign n9539 = ~n9325 & ~n9482;
  assign n9540 = ~n9320 & n9539;
  assign n9541 = n9482 & ~n9485;
  assign n9542 = ~n9540 & ~n9541;
  assign n9543 = ~n9537 & ~n9542;
  assign n9544 = ~n9538 & ~n9543;
  assign n9545 = A430  & A431 ;
  assign n9546 = A430  & ~A431 ;
  assign n9547 = ~A430  & A431 ;
  assign n9548 = ~n9546 & ~n9547;
  assign n9549 = A432  & ~n9548;
  assign n9550 = ~n9545 & ~n9549;
  assign n9551 = A427  & A428 ;
  assign n9552 = A427  & ~A428 ;
  assign n9553 = ~A427  & A428 ;
  assign n9554 = ~n9552 & ~n9553;
  assign n9555 = A429  & ~n9554;
  assign n9556 = ~n9551 & ~n9555;
  assign n9557 = n9550 & ~n9556;
  assign n9558 = ~n9550 & n9556;
  assign n9559 = A429  & ~n9552;
  assign n9560 = ~n9553 & n9559;
  assign n9561 = ~A429  & ~n9554;
  assign n9562 = ~n9560 & ~n9561;
  assign n9563 = A432  & ~n9546;
  assign n9564 = ~n9547 & n9563;
  assign n9565 = ~A432  & ~n9548;
  assign n9566 = ~n9564 & ~n9565;
  assign n9567 = ~n9562 & ~n9566;
  assign n9568 = ~n9558 & n9567;
  assign n9569 = ~n9557 & n9568;
  assign n9570 = ~n9557 & ~n9558;
  assign n9571 = ~n9567 & ~n9570;
  assign n9572 = ~n9569 & ~n9571;
  assign n9573 = ~n9562 & n9566;
  assign n9574 = n9562 & ~n9566;
  assign n9575 = ~n9573 & ~n9574;
  assign n9576 = n9567 & ~n9570;
  assign n9577 = ~n9550 & ~n9556;
  assign n9578 = ~n9576 & ~n9577;
  assign n9579 = ~n9575 & ~n9578;
  assign n9580 = ~n9572 & ~n9579;
  assign n9581 = ~n9572 & ~n9578;
  assign n9582 = A436  & A437 ;
  assign n9583 = A436  & ~A437 ;
  assign n9584 = ~A436  & A437 ;
  assign n9585 = ~n9583 & ~n9584;
  assign n9586 = A438  & ~n9585;
  assign n9587 = ~n9582 & ~n9586;
  assign n9588 = A433  & A434 ;
  assign n9589 = A433  & ~A434 ;
  assign n9590 = ~A433  & A434 ;
  assign n9591 = ~n9589 & ~n9590;
  assign n9592 = A435  & ~n9591;
  assign n9593 = ~n9588 & ~n9592;
  assign n9594 = ~n9587 & n9593;
  assign n9595 = n9587 & ~n9593;
  assign n9596 = ~n9594 & ~n9595;
  assign n9597 = A435  & ~n9589;
  assign n9598 = ~n9590 & n9597;
  assign n9599 = ~A435  & ~n9591;
  assign n9600 = ~n9598 & ~n9599;
  assign n9601 = A438  & ~n9583;
  assign n9602 = ~n9584 & n9601;
  assign n9603 = ~A438  & ~n9585;
  assign n9604 = ~n9602 & ~n9603;
  assign n9605 = ~n9600 & ~n9604;
  assign n9606 = ~n9596 & n9605;
  assign n9607 = ~n9587 & ~n9593;
  assign n9608 = ~n9606 & ~n9607;
  assign n9609 = ~n9594 & n9605;
  assign n9610 = ~n9595 & n9609;
  assign n9611 = ~n9596 & ~n9605;
  assign n9612 = ~n9610 & ~n9611;
  assign n9613 = ~n9608 & ~n9612;
  assign n9614 = ~n9600 & n9604;
  assign n9615 = n9600 & ~n9604;
  assign n9616 = ~n9614 & ~n9615;
  assign n9617 = ~n9575 & ~n9616;
  assign n9618 = ~n9613 & n9617;
  assign n9619 = ~n9581 & n9618;
  assign n9620 = ~n9608 & ~n9616;
  assign n9621 = ~n9612 & ~n9620;
  assign n9622 = ~n9619 & ~n9621;
  assign n9623 = ~n9612 & n9617;
  assign n9624 = ~n9613 & n9623;
  assign n9625 = ~n9581 & ~n9620;
  assign n9626 = n9624 & n9625;
  assign n9627 = ~n9622 & ~n9626;
  assign n9628 = n9580 & ~n9627;
  assign n9629 = ~n9619 & n9621;
  assign n9630 = n9619 & ~n9621;
  assign n9631 = ~n9629 & ~n9630;
  assign n9632 = ~n9580 & ~n9631;
  assign n9633 = ~n9613 & ~n9616;
  assign n9634 = ~n9575 & ~n9581;
  assign n9635 = ~n9633 & n9634;
  assign n9636 = n9633 & ~n9634;
  assign n9637 = ~n9635 & ~n9636;
  assign n9638 = ~A421  & A422 ;
  assign n9639 = A421  & ~A422 ;
  assign n9640 = A423  & ~n9639;
  assign n9641 = ~n9638 & n9640;
  assign n9642 = ~n9638 & ~n9639;
  assign n9643 = ~A423  & ~n9642;
  assign n9644 = ~n9641 & ~n9643;
  assign n9645 = ~A424  & A425 ;
  assign n9646 = A424  & ~A425 ;
  assign n9647 = A426  & ~n9646;
  assign n9648 = ~n9645 & n9647;
  assign n9649 = ~n9645 & ~n9646;
  assign n9650 = ~A426  & ~n9649;
  assign n9651 = ~n9648 & ~n9650;
  assign n9652 = ~n9644 & n9651;
  assign n9653 = n9644 & ~n9651;
  assign n9654 = ~n9652 & ~n9653;
  assign n9655 = A424  & A425 ;
  assign n9656 = A426  & ~n9649;
  assign n9657 = ~n9655 & ~n9656;
  assign n9658 = A421  & A422 ;
  assign n9659 = A423  & ~n9642;
  assign n9660 = ~n9658 & ~n9659;
  assign n9661 = ~n9657 & n9660;
  assign n9662 = n9657 & ~n9660;
  assign n9663 = ~n9661 & ~n9662;
  assign n9664 = ~n9644 & ~n9651;
  assign n9665 = ~n9663 & n9664;
  assign n9666 = ~n9657 & ~n9660;
  assign n9667 = ~n9665 & ~n9666;
  assign n9668 = ~n9661 & n9664;
  assign n9669 = ~n9662 & n9668;
  assign n9670 = ~n9663 & ~n9664;
  assign n9671 = ~n9669 & ~n9670;
  assign n9672 = ~n9667 & ~n9671;
  assign n9673 = ~n9654 & ~n9672;
  assign n9674 = ~A415  & A416 ;
  assign n9675 = A415  & ~A416 ;
  assign n9676 = A417  & ~n9675;
  assign n9677 = ~n9674 & n9676;
  assign n9678 = ~n9674 & ~n9675;
  assign n9679 = ~A417  & ~n9678;
  assign n9680 = ~n9677 & ~n9679;
  assign n9681 = ~A418  & A419 ;
  assign n9682 = A418  & ~A419 ;
  assign n9683 = A420  & ~n9682;
  assign n9684 = ~n9681 & n9683;
  assign n9685 = ~n9681 & ~n9682;
  assign n9686 = ~A420  & ~n9685;
  assign n9687 = ~n9684 & ~n9686;
  assign n9688 = ~n9680 & n9687;
  assign n9689 = n9680 & ~n9687;
  assign n9690 = ~n9688 & ~n9689;
  assign n9691 = A418  & A419 ;
  assign n9692 = A420  & ~n9685;
  assign n9693 = ~n9691 & ~n9692;
  assign n9694 = A415  & A416 ;
  assign n9695 = A417  & ~n9678;
  assign n9696 = ~n9694 & ~n9695;
  assign n9697 = ~n9693 & n9696;
  assign n9698 = n9693 & ~n9696;
  assign n9699 = ~n9697 & ~n9698;
  assign n9700 = ~n9680 & ~n9687;
  assign n9701 = ~n9699 & n9700;
  assign n9702 = ~n9693 & ~n9696;
  assign n9703 = ~n9701 & ~n9702;
  assign n9704 = ~n9697 & n9700;
  assign n9705 = ~n9698 & n9704;
  assign n9706 = ~n9699 & ~n9700;
  assign n9707 = ~n9705 & ~n9706;
  assign n9708 = ~n9703 & ~n9707;
  assign n9709 = ~n9690 & ~n9708;
  assign n9710 = ~n9673 & n9709;
  assign n9711 = n9673 & ~n9709;
  assign n9712 = ~n9710 & ~n9711;
  assign n9713 = ~n9637 & ~n9712;
  assign n9714 = ~n9632 & n9713;
  assign n9715 = ~n9628 & n9714;
  assign n9716 = ~n9628 & ~n9632;
  assign n9717 = ~n9713 & ~n9716;
  assign n9718 = ~n9715 & ~n9717;
  assign n9719 = ~n9690 & ~n9703;
  assign n9720 = ~n9707 & ~n9719;
  assign n9721 = ~n9654 & ~n9690;
  assign n9722 = ~n9672 & n9721;
  assign n9723 = ~n9708 & n9722;
  assign n9724 = ~n9654 & ~n9667;
  assign n9725 = ~n9671 & ~n9724;
  assign n9726 = ~n9723 & n9725;
  assign n9727 = n9723 & ~n9725;
  assign n9728 = ~n9726 & ~n9727;
  assign n9729 = ~n9720 & ~n9728;
  assign n9730 = ~n9723 & ~n9725;
  assign n9731 = ~n9671 & n9721;
  assign n9732 = ~n9672 & n9731;
  assign n9733 = ~n9708 & ~n9724;
  assign n9734 = n9732 & n9733;
  assign n9735 = ~n9730 & ~n9734;
  assign n9736 = n9720 & ~n9735;
  assign n9737 = ~n9729 & ~n9736;
  assign n9738 = ~n9718 & n9737;
  assign n9739 = ~n9632 & ~n9713;
  assign n9740 = ~n9628 & n9739;
  assign n9741 = n9713 & ~n9716;
  assign n9742 = ~n9740 & ~n9741;
  assign n9743 = ~n9737 & ~n9742;
  assign n9744 = ~n9738 & ~n9743;
  assign n9745 = A442  & A443 ;
  assign n9746 = A442  & ~A443 ;
  assign n9747 = ~A442  & A443 ;
  assign n9748 = ~n9746 & ~n9747;
  assign n9749 = A444  & ~n9748;
  assign n9750 = ~n9745 & ~n9749;
  assign n9751 = A439  & A440 ;
  assign n9752 = A439  & ~A440 ;
  assign n9753 = ~A439  & A440 ;
  assign n9754 = ~n9752 & ~n9753;
  assign n9755 = A441  & ~n9754;
  assign n9756 = ~n9751 & ~n9755;
  assign n9757 = n9750 & ~n9756;
  assign n9758 = ~n9750 & n9756;
  assign n9759 = A441  & ~n9752;
  assign n9760 = ~n9753 & n9759;
  assign n9761 = ~A441  & ~n9754;
  assign n9762 = ~n9760 & ~n9761;
  assign n9763 = A444  & ~n9746;
  assign n9764 = ~n9747 & n9763;
  assign n9765 = ~A444  & ~n9748;
  assign n9766 = ~n9764 & ~n9765;
  assign n9767 = ~n9762 & ~n9766;
  assign n9768 = ~n9758 & n9767;
  assign n9769 = ~n9757 & n9768;
  assign n9770 = ~n9757 & ~n9758;
  assign n9771 = ~n9767 & ~n9770;
  assign n9772 = ~n9769 & ~n9771;
  assign n9773 = ~n9762 & n9766;
  assign n9774 = n9762 & ~n9766;
  assign n9775 = ~n9773 & ~n9774;
  assign n9776 = n9767 & ~n9770;
  assign n9777 = ~n9750 & ~n9756;
  assign n9778 = ~n9776 & ~n9777;
  assign n9779 = ~n9775 & ~n9778;
  assign n9780 = ~n9772 & ~n9779;
  assign n9781 = ~n9772 & ~n9778;
  assign n9782 = A448  & A449 ;
  assign n9783 = A448  & ~A449 ;
  assign n9784 = ~A448  & A449 ;
  assign n9785 = ~n9783 & ~n9784;
  assign n9786 = A450  & ~n9785;
  assign n9787 = ~n9782 & ~n9786;
  assign n9788 = A445  & A446 ;
  assign n9789 = A445  & ~A446 ;
  assign n9790 = ~A445  & A446 ;
  assign n9791 = ~n9789 & ~n9790;
  assign n9792 = A447  & ~n9791;
  assign n9793 = ~n9788 & ~n9792;
  assign n9794 = ~n9787 & n9793;
  assign n9795 = n9787 & ~n9793;
  assign n9796 = ~n9794 & ~n9795;
  assign n9797 = A447  & ~n9789;
  assign n9798 = ~n9790 & n9797;
  assign n9799 = ~A447  & ~n9791;
  assign n9800 = ~n9798 & ~n9799;
  assign n9801 = A450  & ~n9783;
  assign n9802 = ~n9784 & n9801;
  assign n9803 = ~A450  & ~n9785;
  assign n9804 = ~n9802 & ~n9803;
  assign n9805 = ~n9800 & ~n9804;
  assign n9806 = ~n9796 & n9805;
  assign n9807 = ~n9787 & ~n9793;
  assign n9808 = ~n9806 & ~n9807;
  assign n9809 = ~n9794 & n9805;
  assign n9810 = ~n9795 & n9809;
  assign n9811 = ~n9796 & ~n9805;
  assign n9812 = ~n9810 & ~n9811;
  assign n9813 = ~n9808 & ~n9812;
  assign n9814 = ~n9800 & n9804;
  assign n9815 = n9800 & ~n9804;
  assign n9816 = ~n9814 & ~n9815;
  assign n9817 = ~n9775 & ~n9816;
  assign n9818 = ~n9813 & n9817;
  assign n9819 = ~n9781 & n9818;
  assign n9820 = ~n9808 & ~n9816;
  assign n9821 = ~n9812 & ~n9820;
  assign n9822 = ~n9819 & n9821;
  assign n9823 = n9819 & ~n9821;
  assign n9824 = ~n9822 & ~n9823;
  assign n9825 = ~n9780 & ~n9824;
  assign n9826 = ~n9819 & ~n9821;
  assign n9827 = ~n9812 & n9817;
  assign n9828 = ~n9813 & n9827;
  assign n9829 = ~n9781 & ~n9820;
  assign n9830 = n9828 & n9829;
  assign n9831 = ~n9826 & ~n9830;
  assign n9832 = n9780 & ~n9831;
  assign n9833 = ~n9825 & ~n9832;
  assign n9834 = A454  & A455 ;
  assign n9835 = A454  & ~A455 ;
  assign n9836 = ~A454  & A455 ;
  assign n9837 = ~n9835 & ~n9836;
  assign n9838 = A456  & ~n9837;
  assign n9839 = ~n9834 & ~n9838;
  assign n9840 = A451  & A452 ;
  assign n9841 = A451  & ~A452 ;
  assign n9842 = ~A451  & A452 ;
  assign n9843 = ~n9841 & ~n9842;
  assign n9844 = A453  & ~n9843;
  assign n9845 = ~n9840 & ~n9844;
  assign n9846 = n9839 & ~n9845;
  assign n9847 = ~n9839 & n9845;
  assign n9848 = A453  & ~n9841;
  assign n9849 = ~n9842 & n9848;
  assign n9850 = ~A453  & ~n9843;
  assign n9851 = ~n9849 & ~n9850;
  assign n9852 = A456  & ~n9835;
  assign n9853 = ~n9836 & n9852;
  assign n9854 = ~A456  & ~n9837;
  assign n9855 = ~n9853 & ~n9854;
  assign n9856 = ~n9851 & ~n9855;
  assign n9857 = ~n9847 & n9856;
  assign n9858 = ~n9846 & n9857;
  assign n9859 = ~n9846 & ~n9847;
  assign n9860 = ~n9856 & ~n9859;
  assign n9861 = ~n9858 & ~n9860;
  assign n9862 = ~n9851 & n9855;
  assign n9863 = n9851 & ~n9855;
  assign n9864 = ~n9862 & ~n9863;
  assign n9865 = n9856 & ~n9859;
  assign n9866 = ~n9839 & ~n9845;
  assign n9867 = ~n9865 & ~n9866;
  assign n9868 = ~n9864 & ~n9867;
  assign n9869 = ~n9861 & ~n9868;
  assign n9870 = ~n9861 & ~n9867;
  assign n9871 = A460  & A461 ;
  assign n9872 = A460  & ~A461 ;
  assign n9873 = ~A460  & A461 ;
  assign n9874 = ~n9872 & ~n9873;
  assign n9875 = A462  & ~n9874;
  assign n9876 = ~n9871 & ~n9875;
  assign n9877 = A457  & A458 ;
  assign n9878 = A457  & ~A458 ;
  assign n9879 = ~A457  & A458 ;
  assign n9880 = ~n9878 & ~n9879;
  assign n9881 = A459  & ~n9880;
  assign n9882 = ~n9877 & ~n9881;
  assign n9883 = ~n9876 & n9882;
  assign n9884 = n9876 & ~n9882;
  assign n9885 = ~n9883 & ~n9884;
  assign n9886 = A459  & ~n9878;
  assign n9887 = ~n9879 & n9886;
  assign n9888 = ~A459  & ~n9880;
  assign n9889 = ~n9887 & ~n9888;
  assign n9890 = A462  & ~n9872;
  assign n9891 = ~n9873 & n9890;
  assign n9892 = ~A462  & ~n9874;
  assign n9893 = ~n9891 & ~n9892;
  assign n9894 = ~n9889 & ~n9893;
  assign n9895 = ~n9885 & n9894;
  assign n9896 = ~n9876 & ~n9882;
  assign n9897 = ~n9895 & ~n9896;
  assign n9898 = ~n9883 & n9894;
  assign n9899 = ~n9884 & n9898;
  assign n9900 = ~n9885 & ~n9894;
  assign n9901 = ~n9899 & ~n9900;
  assign n9902 = ~n9897 & ~n9901;
  assign n9903 = ~n9889 & n9893;
  assign n9904 = n9889 & ~n9893;
  assign n9905 = ~n9903 & ~n9904;
  assign n9906 = ~n9864 & ~n9905;
  assign n9907 = ~n9902 & n9906;
  assign n9908 = ~n9870 & n9907;
  assign n9909 = ~n9897 & ~n9905;
  assign n9910 = ~n9901 & ~n9909;
  assign n9911 = ~n9908 & ~n9910;
  assign n9912 = ~n9901 & n9906;
  assign n9913 = ~n9902 & n9912;
  assign n9914 = ~n9870 & ~n9909;
  assign n9915 = n9913 & n9914;
  assign n9916 = ~n9911 & ~n9915;
  assign n9917 = n9869 & ~n9916;
  assign n9918 = ~n9908 & n9910;
  assign n9919 = n9908 & ~n9910;
  assign n9920 = ~n9918 & ~n9919;
  assign n9921 = ~n9869 & ~n9920;
  assign n9922 = ~n9902 & ~n9905;
  assign n9923 = ~n9864 & ~n9870;
  assign n9924 = ~n9922 & n9923;
  assign n9925 = n9922 & ~n9923;
  assign n9926 = ~n9924 & ~n9925;
  assign n9927 = ~n9813 & ~n9816;
  assign n9928 = ~n9775 & ~n9781;
  assign n9929 = ~n9927 & n9928;
  assign n9930 = n9927 & ~n9928;
  assign n9931 = ~n9929 & ~n9930;
  assign n9932 = ~n9926 & ~n9931;
  assign n9933 = ~n9921 & ~n9932;
  assign n9934 = ~n9917 & n9933;
  assign n9935 = ~n9917 & ~n9921;
  assign n9936 = n9932 & ~n9935;
  assign n9937 = ~n9934 & ~n9936;
  assign n9938 = ~n9833 & ~n9937;
  assign n9939 = ~n9921 & n9932;
  assign n9940 = ~n9917 & n9939;
  assign n9941 = ~n9932 & ~n9935;
  assign n9942 = ~n9940 & ~n9941;
  assign n9943 = n9833 & ~n9942;
  assign n9944 = ~n9926 & n9931;
  assign n9945 = n9926 & ~n9931;
  assign n9946 = ~n9944 & ~n9945;
  assign n9947 = ~n9637 & n9712;
  assign n9948 = n9637 & ~n9712;
  assign n9949 = ~n9947 & ~n9948;
  assign n9950 = ~n9946 & ~n9949;
  assign n9951 = ~n9943 & ~n9950;
  assign n9952 = ~n9938 & n9951;
  assign n9953 = ~n9938 & ~n9943;
  assign n9954 = n9950 & ~n9953;
  assign n9955 = ~n9952 & ~n9954;
  assign n9956 = ~n9744 & ~n9955;
  assign n9957 = ~n9943 & n9950;
  assign n9958 = ~n9938 & n9957;
  assign n9959 = ~n9950 & ~n9953;
  assign n9960 = ~n9958 & ~n9959;
  assign n9961 = n9744 & ~n9960;
  assign n9962 = ~n9946 & n9949;
  assign n9963 = n9946 & ~n9949;
  assign n9964 = ~n9962 & ~n9963;
  assign n9965 = ~n9328 & n9481;
  assign n9966 = n9328 & ~n9481;
  assign n9967 = ~n9965 & ~n9966;
  assign n9968 = ~n9964 & ~n9967;
  assign n9969 = ~n9961 & ~n9968;
  assign n9970 = ~n9956 & n9969;
  assign n9971 = ~n9956 & ~n9961;
  assign n9972 = n9968 & ~n9971;
  assign n9973 = ~n9970 & ~n9972;
  assign n9974 = ~n9544 & ~n9973;
  assign n9975 = ~n9961 & n9968;
  assign n9976 = ~n9956 & n9975;
  assign n9977 = ~n9968 & ~n9971;
  assign n9978 = ~n9976 & ~n9977;
  assign n9979 = n9544 & ~n9978;
  assign n9980 = ~n9964 & n9967;
  assign n9981 = n9964 & ~n9967;
  assign n9982 = ~n9980 & ~n9981;
  assign n9983 = ~n8692 & n9001;
  assign n9984 = n8692 & ~n9001;
  assign n9985 = ~n9983 & ~n9984;
  assign n9986 = ~n9982 & ~n9985;
  assign n9987 = ~n9979 & ~n9986;
  assign n9988 = ~n9974 & n9987;
  assign n9989 = ~n9974 & ~n9979;
  assign n9990 = n9986 & ~n9989;
  assign n9991 = ~n9988 & ~n9990;
  assign n9992 = ~n9126 & ~n9991;
  assign n9993 = ~n9979 & n9986;
  assign n9994 = ~n9974 & n9993;
  assign n9995 = ~n9986 & ~n9989;
  assign n9996 = ~n9994 & ~n9995;
  assign n9997 = n9126 & ~n9996;
  assign n9998 = ~n9982 & n9985;
  assign n9999 = n9982 & ~n9985;
  assign n10000 = ~n9998 & ~n9999;
  assign n10001 = ~n7402 & n8023;
  assign n10002 = n7402 & ~n8023;
  assign n10003 = ~n10001 & ~n10002;
  assign n10004 = ~n10000 & ~n10003;
  assign n10005 = ~n9997 & ~n10004;
  assign n10006 = ~n9992 & n10005;
  assign n10007 = ~n9992 & ~n9997;
  assign n10008 = n10004 & ~n10007;
  assign n10009 = ~n10006 & ~n10008;
  assign n10010 = ~n8272 & ~n10009;
  assign n10011 = ~n9997 & n10004;
  assign n10012 = ~n9992 & n10011;
  assign n10013 = ~n10004 & ~n10007;
  assign n10014 = ~n10012 & ~n10013;
  assign n10015 = n8272 & ~n10014;
  assign n10016 = ~n10000 & n10003;
  assign n10017 = n10000 & ~n10003;
  assign n10018 = ~n10016 & ~n10017;
  assign n10019 = ~n5676 & n6297;
  assign n10020 = ~n5673 & ~n6297;
  assign n10021 = ~n5675 & n10020;
  assign n10022 = ~n10019 & ~n10021;
  assign n10023 = ~n10018 & ~n10022;
  assign n10024 = ~n10015 & ~n10023;
  assign n10025 = ~n10010 & n10024;
  assign n10026 = ~n10010 & ~n10015;
  assign n10027 = n10023 & ~n10026;
  assign n10028 = ~n10025 & ~n10027;
  assign n10029 = ~n6546 & ~n10028;
  assign n10030 = ~n3972 & n3975;
  assign n10031 = n3972 & ~n3975;
  assign n10032 = ~n10030 & ~n10031;
  assign n10033 = ~n10018 & n10022;
  assign n10034 = n10018 & ~n10022;
  assign n10035 = ~n10033 & ~n10034;
  assign n10036 = ~n10032 & ~n10035;
  assign n10037 = ~n10015 & n10023;
  assign n10038 = ~n10010 & n10037;
  assign n10039 = ~n10023 & ~n10026;
  assign n10040 = ~n10038 & ~n10039;
  assign n10041 = n6546 & ~n10040;
  assign n10042 = ~n10036 & ~n10041;
  assign n10043 = ~n10029 & n10042;
  assign n10044 = ~n4472 & ~n10043;
  assign n10045 = ~n10029 & ~n10041;
  assign n10046 = n10036 & ~n10045;
  assign n10047 = ~n10044 & ~n10046;
  assign n10048 = ~n6546 & ~n10025;
  assign n10049 = ~n10027 & ~n10048;
  assign n10050 = ~n6539 & ~n6542;
  assign n10051 = ~n6543 & ~n10050;
  assign n10052 = ~n4890 & ~n5663;
  assign n10053 = ~n5665 & ~n10052;
  assign n10054 = ~n5218 & ~n5645;
  assign n10055 = ~n5647 & ~n10054;
  assign n10056 = ~n5211 & ~n5214;
  assign n10057 = ~n5215 & ~n10056;
  assign n10058 = n5172 & ~n5207;
  assign n10059 = ~n5208 & ~n10058;
  assign n10060 = ~n5193 & ~n5194;
  assign n10061 = ~n5190 & ~n10060;
  assign n10062 = ~n5177 & ~n5180;
  assign n10063 = ~n5187 & ~n10062;
  assign n10064 = ~n10061 & n10063;
  assign n10065 = ~n5190 & ~n10063;
  assign n10066 = ~n10060 & n10065;
  assign n10067 = ~n5109 & ~n5126;
  assign n10068 = ~n5122 & ~n10067;
  assign n10069 = ~n10066 & n10068;
  assign n10070 = ~n10064 & n10069;
  assign n10071 = ~n10064 & ~n10066;
  assign n10072 = ~n10068 & ~n10071;
  assign n10073 = ~n10070 & ~n10072;
  assign n10074 = ~n10059 & ~n10073;
  assign n10075 = ~n5208 & ~n10070;
  assign n10076 = ~n10058 & n10075;
  assign n10077 = ~n10072 & n10076;
  assign n10078 = ~n10074 & ~n10077;
  assign n10079 = ~n4979 & ~n5080;
  assign n10080 = ~n5082 & ~n10079;
  assign n10081 = n4926 & ~n4972;
  assign n10082 = ~n4976 & ~n10081;
  assign n10083 = ~n4958 & ~n4962;
  assign n10084 = ~n4954 & ~n10083;
  assign n10085 = ~n4918 & ~n4921;
  assign n10086 = ~n4924 & ~n10085;
  assign n10087 = ~n10084 & n10086;
  assign n10088 = n10084 & ~n10086;
  assign n10089 = ~n10087 & ~n10088;
  assign n10090 = ~n10082 & ~n10089;
  assign n10091 = ~n4976 & ~n10087;
  assign n10092 = ~n10088 & n10091;
  assign n10093 = ~n10081 & n10092;
  assign n10094 = ~n10090 & ~n10093;
  assign n10095 = n5015 & ~n5057;
  assign n10096 = ~n5061 & ~n10095;
  assign n10097 = ~n5047 & ~n5051;
  assign n10098 = ~n5043 & ~n10097;
  assign n10099 = ~n5007 & ~n5010;
  assign n10100 = ~n5013 & ~n10099;
  assign n10101 = ~n10098 & n10100;
  assign n10102 = n10098 & ~n10100;
  assign n10103 = ~n10101 & ~n10102;
  assign n10104 = ~n10096 & ~n10103;
  assign n10105 = ~n5061 & ~n10101;
  assign n10106 = ~n10102 & n10105;
  assign n10107 = ~n10095 & n10106;
  assign n10108 = ~n10104 & ~n10107;
  assign n10109 = ~n10094 & n10108;
  assign n10110 = n10094 & ~n10108;
  assign n10111 = ~n10109 & ~n10110;
  assign n10112 = ~n10080 & ~n10111;
  assign n10113 = n10080 & n10111;
  assign n10114 = ~n10112 & ~n10113;
  assign n10115 = ~n10078 & n10114;
  assign n10116 = n10078 & ~n10114;
  assign n10117 = ~n10115 & ~n10116;
  assign n10118 = ~n10057 & ~n10117;
  assign n10119 = n10057 & n10117;
  assign n10120 = ~n10118 & ~n10119;
  assign n10121 = ~n5418 & ~n5626;
  assign n10122 = ~n5628 & ~n10121;
  assign n10123 = ~n5411 & ~n5414;
  assign n10124 = ~n5415 & ~n10123;
  assign n10125 = n5394 & ~n5404;
  assign n10126 = ~n5408 & ~n10125;
  assign n10127 = ~n5328 & ~n5345;
  assign n10128 = ~n5341 & ~n10127;
  assign n10129 = ~n5364 & ~n5381;
  assign n10130 = ~n5377 & ~n10129;
  assign n10131 = ~n10128 & n10130;
  assign n10132 = n10128 & ~n10130;
  assign n10133 = ~n10131 & ~n10132;
  assign n10134 = ~n10126 & ~n10133;
  assign n10135 = ~n5408 & ~n10131;
  assign n10136 = ~n10132 & n10135;
  assign n10137 = ~n10125 & n10136;
  assign n10138 = ~n10134 & ~n10137;
  assign n10139 = n5254 & ~n5296;
  assign n10140 = ~n5300 & ~n10139;
  assign n10141 = ~n5286 & ~n5290;
  assign n10142 = ~n5282 & ~n10141;
  assign n10143 = ~n5246 & ~n5249;
  assign n10144 = ~n5252 & ~n10143;
  assign n10145 = ~n10142 & n10144;
  assign n10146 = n10142 & ~n10144;
  assign n10147 = ~n10145 & ~n10146;
  assign n10148 = ~n10140 & ~n10147;
  assign n10149 = ~n5300 & ~n10145;
  assign n10150 = ~n10146 & n10149;
  assign n10151 = ~n10139 & n10150;
  assign n10152 = ~n10148 & ~n10151;
  assign n10153 = ~n10138 & n10152;
  assign n10154 = n10138 & ~n10152;
  assign n10155 = ~n10153 & ~n10154;
  assign n10156 = ~n10124 & ~n10155;
  assign n10157 = n10124 & n10155;
  assign n10158 = ~n10156 & ~n10157;
  assign n10159 = ~n5507 & ~n5608;
  assign n10160 = ~n5610 & ~n10159;
  assign n10161 = n5454 & ~n5500;
  assign n10162 = ~n5504 & ~n10161;
  assign n10163 = ~n5486 & ~n5490;
  assign n10164 = ~n5482 & ~n10163;
  assign n10165 = ~n5446 & ~n5449;
  assign n10166 = ~n5452 & ~n10165;
  assign n10167 = ~n10164 & n10166;
  assign n10168 = n10164 & ~n10166;
  assign n10169 = ~n10167 & ~n10168;
  assign n10170 = ~n10162 & ~n10169;
  assign n10171 = ~n5504 & ~n10167;
  assign n10172 = ~n10168 & n10171;
  assign n10173 = ~n10161 & n10172;
  assign n10174 = ~n10170 & ~n10173;
  assign n10175 = n5543 & ~n5585;
  assign n10176 = ~n5589 & ~n10175;
  assign n10177 = ~n5575 & ~n5579;
  assign n10178 = ~n5571 & ~n10177;
  assign n10179 = ~n5535 & ~n5538;
  assign n10180 = ~n5541 & ~n10179;
  assign n10181 = ~n10178 & n10180;
  assign n10182 = n10178 & ~n10180;
  assign n10183 = ~n10181 & ~n10182;
  assign n10184 = ~n10176 & ~n10183;
  assign n10185 = ~n5589 & ~n10181;
  assign n10186 = ~n10182 & n10185;
  assign n10187 = ~n10175 & n10186;
  assign n10188 = ~n10184 & ~n10187;
  assign n10189 = ~n10174 & n10188;
  assign n10190 = n10174 & ~n10188;
  assign n10191 = ~n10189 & ~n10190;
  assign n10192 = ~n10160 & ~n10191;
  assign n10193 = n10160 & n10191;
  assign n10194 = ~n10192 & ~n10193;
  assign n10195 = ~n10158 & n10194;
  assign n10196 = n10158 & ~n10194;
  assign n10197 = ~n10195 & ~n10196;
  assign n10198 = ~n10122 & ~n10197;
  assign n10199 = n10122 & n10197;
  assign n10200 = ~n10198 & ~n10199;
  assign n10201 = ~n10120 & n10200;
  assign n10202 = n10120 & ~n10200;
  assign n10203 = ~n10201 & ~n10202;
  assign n10204 = n10055 & n10203;
  assign n10205 = ~n10055 & ~n10203;
  assign n10206 = ~n4883 & ~n4886;
  assign n10207 = ~n4887 & ~n10206;
  assign n10208 = ~n4876 & ~n4879;
  assign n10209 = ~n4880 & ~n10208;
  assign n10210 = n4859 & ~n4869;
  assign n10211 = ~n4873 & ~n10210;
  assign n10212 = ~n4766 & ~n4783;
  assign n10213 = ~n4779 & ~n10212;
  assign n10214 = ~n4802 & ~n4819;
  assign n10215 = ~n4815 & ~n10214;
  assign n10216 = ~n10213 & n10215;
  assign n10217 = n10213 & ~n10215;
  assign n10218 = ~n10216 & ~n10217;
  assign n10219 = ~n10211 & ~n10218;
  assign n10220 = ~n4873 & ~n10216;
  assign n10221 = ~n10217 & n10220;
  assign n10222 = ~n10210 & n10221;
  assign n10223 = ~n10219 & ~n10222;
  assign n10224 = n4835 & ~n4841;
  assign n10225 = ~n4845 & ~n10224;
  assign n10226 = ~n4691 & ~n4708;
  assign n10227 = ~n4704 & ~n10226;
  assign n10228 = ~n4727 & ~n4744;
  assign n10229 = ~n4740 & ~n10228;
  assign n10230 = ~n10227 & n10229;
  assign n10231 = n10227 & ~n10229;
  assign n10232 = ~n10230 & ~n10231;
  assign n10233 = ~n10225 & ~n10232;
  assign n10234 = ~n4845 & ~n10230;
  assign n10235 = ~n10231 & n10234;
  assign n10236 = ~n10224 & n10235;
  assign n10237 = ~n10233 & ~n10236;
  assign n10238 = ~n10223 & n10237;
  assign n10239 = n10223 & ~n10237;
  assign n10240 = ~n10238 & ~n10239;
  assign n10241 = ~n10209 & ~n10240;
  assign n10242 = n10209 & n10240;
  assign n10243 = ~n10241 & ~n10242;
  assign n10244 = ~n4561 & ~n4662;
  assign n10245 = ~n4664 & ~n10244;
  assign n10246 = n4508 & ~n4554;
  assign n10247 = ~n4558 & ~n10246;
  assign n10248 = ~n4540 & ~n4544;
  assign n10249 = ~n4536 & ~n10248;
  assign n10250 = ~n4500 & ~n4503;
  assign n10251 = ~n4506 & ~n10250;
  assign n10252 = ~n10249 & n10251;
  assign n10253 = n10249 & ~n10251;
  assign n10254 = ~n10252 & ~n10253;
  assign n10255 = ~n10247 & ~n10254;
  assign n10256 = ~n4558 & ~n10252;
  assign n10257 = ~n10253 & n10256;
  assign n10258 = ~n10246 & n10257;
  assign n10259 = ~n10255 & ~n10258;
  assign n10260 = n4597 & ~n4639;
  assign n10261 = ~n4643 & ~n10260;
  assign n10262 = ~n4629 & ~n4633;
  assign n10263 = ~n4625 & ~n10262;
  assign n10264 = ~n4589 & ~n4592;
  assign n10265 = ~n4595 & ~n10264;
  assign n10266 = ~n10263 & n10265;
  assign n10267 = n10263 & ~n10265;
  assign n10268 = ~n10266 & ~n10267;
  assign n10269 = ~n10261 & ~n10268;
  assign n10270 = ~n4643 & ~n10266;
  assign n10271 = ~n10267 & n10270;
  assign n10272 = ~n10260 & n10271;
  assign n10273 = ~n10269 & ~n10272;
  assign n10274 = ~n10259 & n10273;
  assign n10275 = n10259 & ~n10273;
  assign n10276 = ~n10274 & ~n10275;
  assign n10277 = ~n10245 & ~n10276;
  assign n10278 = n10245 & n10276;
  assign n10279 = ~n10277 & ~n10278;
  assign n10280 = ~n10243 & n10279;
  assign n10281 = n10243 & ~n10279;
  assign n10282 = ~n10280 & ~n10281;
  assign n10283 = ~n10207 & ~n10282;
  assign n10284 = n10207 & n10282;
  assign n10285 = ~n10283 & ~n10284;
  assign n10286 = ~n10205 & ~n10285;
  assign n10287 = ~n10204 & n10286;
  assign n10288 = ~n10204 & ~n10205;
  assign n10289 = n10285 & ~n10288;
  assign n10290 = ~n10287 & ~n10289;
  assign n10291 = n10053 & n10290;
  assign n10292 = ~n10053 & ~n10290;
  assign n10293 = ~n6532 & ~n6535;
  assign n10294 = ~n6536 & ~n10293;
  assign n10295 = ~n6525 & ~n6528;
  assign n10296 = ~n6529 & ~n10295;
  assign n10297 = ~n6518 & ~n6521;
  assign n10298 = ~n6522 & ~n10297;
  assign n10299 = n6501 & ~n6511;
  assign n10300 = ~n6515 & ~n10299;
  assign n10301 = ~n6230 & ~n6247;
  assign n10302 = ~n6243 & ~n10301;
  assign n10303 = ~n6266 & ~n6283;
  assign n10304 = ~n6279 & ~n10303;
  assign n10305 = ~n10302 & n10304;
  assign n10306 = n10302 & ~n10304;
  assign n10307 = ~n10305 & ~n10306;
  assign n10308 = ~n10300 & ~n10307;
  assign n10309 = ~n6515 & ~n10305;
  assign n10310 = ~n10306 & n10309;
  assign n10311 = ~n10299 & n10310;
  assign n10312 = ~n10308 & ~n10311;
  assign n10313 = n6477 & ~n6483;
  assign n10314 = ~n6487 & ~n10313;
  assign n10315 = ~n6155 & ~n6172;
  assign n10316 = ~n6168 & ~n10315;
  assign n10317 = ~n6191 & ~n6208;
  assign n10318 = ~n6204 & ~n10317;
  assign n10319 = ~n10316 & n10318;
  assign n10320 = n10316 & ~n10318;
  assign n10321 = ~n10319 & ~n10320;
  assign n10322 = ~n10314 & ~n10321;
  assign n10323 = ~n6487 & ~n10319;
  assign n10324 = ~n10320 & n10323;
  assign n10325 = ~n10313 & n10324;
  assign n10326 = ~n10322 & ~n10325;
  assign n10327 = ~n10312 & n10326;
  assign n10328 = n10312 & ~n10326;
  assign n10329 = ~n10327 & ~n10328;
  assign n10330 = ~n10298 & ~n10329;
  assign n10331 = n10298 & n10329;
  assign n10332 = ~n10330 & ~n10331;
  assign n10333 = ~n6439 & ~n6460;
  assign n10334 = ~n6462 & ~n10333;
  assign n10335 = n6422 & ~n6432;
  assign n10336 = ~n6436 & ~n10335;
  assign n10337 = ~n6077 & ~n6094;
  assign n10338 = ~n6090 & ~n10337;
  assign n10339 = ~n6113 & ~n6130;
  assign n10340 = ~n6126 & ~n10339;
  assign n10341 = ~n10338 & n10340;
  assign n10342 = n10338 & ~n10340;
  assign n10343 = ~n10341 & ~n10342;
  assign n10344 = ~n10336 & ~n10343;
  assign n10345 = ~n6436 & ~n10341;
  assign n10346 = ~n10342 & n10345;
  assign n10347 = ~n10335 & n10346;
  assign n10348 = ~n10344 & ~n10347;
  assign n10349 = n6441 & ~n6447;
  assign n10350 = ~n6451 & ~n10349;
  assign n10351 = ~n6002 & ~n6019;
  assign n10352 = ~n6015 & ~n10351;
  assign n10353 = ~n6038 & ~n6055;
  assign n10354 = ~n6051 & ~n10353;
  assign n10355 = ~n10352 & n10354;
  assign n10356 = n10352 & ~n10354;
  assign n10357 = ~n10355 & ~n10356;
  assign n10358 = ~n10350 & ~n10357;
  assign n10359 = ~n6451 & ~n10355;
  assign n10360 = ~n10356 & n10359;
  assign n10361 = ~n10349 & n10360;
  assign n10362 = ~n10358 & ~n10361;
  assign n10363 = ~n10348 & n10362;
  assign n10364 = n10348 & ~n10362;
  assign n10365 = ~n10363 & ~n10364;
  assign n10366 = ~n10334 & ~n10365;
  assign n10367 = n10334 & n10365;
  assign n10368 = ~n10366 & ~n10367;
  assign n10369 = ~n10332 & n10368;
  assign n10370 = n10332 & ~n10368;
  assign n10371 = ~n10369 & ~n10370;
  assign n10372 = ~n10296 & ~n10371;
  assign n10373 = n10296 & n10371;
  assign n10374 = ~n10372 & ~n10373;
  assign n10375 = ~n6353 & ~n6405;
  assign n10376 = ~n6407 & ~n10375;
  assign n10377 = ~n6346 & ~n6349;
  assign n10378 = ~n6350 & ~n10377;
  assign n10379 = n6329 & ~n6339;
  assign n10380 = ~n6343 & ~n10379;
  assign n10381 = ~n5921 & ~n5938;
  assign n10382 = ~n5934 & ~n10381;
  assign n10383 = ~n5957 & ~n5974;
  assign n10384 = ~n5970 & ~n10383;
  assign n10385 = ~n10382 & n10384;
  assign n10386 = n10382 & ~n10384;
  assign n10387 = ~n10385 & ~n10386;
  assign n10388 = ~n10380 & ~n10387;
  assign n10389 = ~n6343 & ~n10385;
  assign n10390 = ~n10386 & n10389;
  assign n10391 = ~n10379 & n10390;
  assign n10392 = ~n10388 & ~n10391;
  assign n10393 = n6305 & ~n6311;
  assign n10394 = ~n6315 & ~n10393;
  assign n10395 = ~n5846 & ~n5863;
  assign n10396 = ~n5859 & ~n10395;
  assign n10397 = ~n5882 & ~n5899;
  assign n10398 = ~n5895 & ~n10397;
  assign n10399 = ~n10396 & n10398;
  assign n10400 = n10396 & ~n10398;
  assign n10401 = ~n10399 & ~n10400;
  assign n10402 = ~n10394 & ~n10401;
  assign n10403 = ~n6315 & ~n10399;
  assign n10404 = ~n10400 & n10403;
  assign n10405 = ~n10393 & n10404;
  assign n10406 = ~n10402 & ~n10405;
  assign n10407 = ~n10392 & n10406;
  assign n10408 = n10392 & ~n10406;
  assign n10409 = ~n10407 & ~n10408;
  assign n10410 = ~n10378 & ~n10409;
  assign n10411 = n10378 & n10409;
  assign n10412 = ~n10410 & ~n10411;
  assign n10413 = ~n6372 & ~n6393;
  assign n10414 = ~n6395 & ~n10413;
  assign n10415 = n6355 & ~n6365;
  assign n10416 = ~n6369 & ~n10415;
  assign n10417 = ~n5768 & ~n5785;
  assign n10418 = ~n5781 & ~n10417;
  assign n10419 = ~n5804 & ~n5821;
  assign n10420 = ~n5817 & ~n10419;
  assign n10421 = ~n10418 & n10420;
  assign n10422 = n10418 & ~n10420;
  assign n10423 = ~n10421 & ~n10422;
  assign n10424 = ~n10416 & ~n10423;
  assign n10425 = ~n6369 & ~n10421;
  assign n10426 = ~n10422 & n10425;
  assign n10427 = ~n10415 & n10426;
  assign n10428 = ~n10424 & ~n10427;
  assign n10429 = n6374 & ~n6380;
  assign n10430 = ~n6384 & ~n10429;
  assign n10431 = ~n5693 & ~n5710;
  assign n10432 = ~n5706 & ~n10431;
  assign n10433 = ~n5729 & ~n5746;
  assign n10434 = ~n5742 & ~n10433;
  assign n10435 = ~n10432 & n10434;
  assign n10436 = n10432 & ~n10434;
  assign n10437 = ~n10435 & ~n10436;
  assign n10438 = ~n10430 & ~n10437;
  assign n10439 = ~n6384 & ~n10435;
  assign n10440 = ~n10436 & n10439;
  assign n10441 = ~n10429 & n10440;
  assign n10442 = ~n10438 & ~n10441;
  assign n10443 = ~n10428 & n10442;
  assign n10444 = n10428 & ~n10442;
  assign n10445 = ~n10443 & ~n10444;
  assign n10446 = ~n10414 & ~n10445;
  assign n10447 = n10414 & n10445;
  assign n10448 = ~n10446 & ~n10447;
  assign n10449 = ~n10412 & n10448;
  assign n10450 = n10412 & ~n10448;
  assign n10451 = ~n10449 & ~n10450;
  assign n10452 = ~n10376 & ~n10451;
  assign n10453 = n10376 & n10451;
  assign n10454 = ~n10452 & ~n10453;
  assign n10455 = ~n10374 & n10454;
  assign n10456 = n10374 & ~n10454;
  assign n10457 = ~n10455 & ~n10456;
  assign n10458 = ~n10294 & ~n10457;
  assign n10459 = n10294 & n10457;
  assign n10460 = ~n10458 & ~n10459;
  assign n10461 = ~n10292 & ~n10460;
  assign n10462 = ~n10291 & n10461;
  assign n10463 = ~n10291 & ~n10292;
  assign n10464 = n10460 & ~n10463;
  assign n10465 = ~n10462 & ~n10464;
  assign n10466 = ~n10051 & ~n10465;
  assign n10467 = n10051 & n10465;
  assign n10468 = ~n10466 & ~n10467;
  assign n10469 = ~n8272 & ~n10006;
  assign n10470 = ~n10008 & ~n10469;
  assign n10471 = ~n8265 & ~n8268;
  assign n10472 = ~n8269 & ~n10471;
  assign n10473 = ~n8258 & ~n8261;
  assign n10474 = ~n8262 & ~n10473;
  assign n10475 = ~n8251 & ~n8254;
  assign n10476 = ~n8255 & ~n10475;
  assign n10477 = ~n8244 & ~n8247;
  assign n10478 = ~n8248 & ~n10477;
  assign n10479 = n8227 & ~n8237;
  assign n10480 = ~n8241 & ~n10479;
  assign n10481 = ~n7956 & ~n7973;
  assign n10482 = ~n7969 & ~n10481;
  assign n10483 = ~n7992 & ~n8009;
  assign n10484 = ~n8005 & ~n10483;
  assign n10485 = ~n10482 & n10484;
  assign n10486 = n10482 & ~n10484;
  assign n10487 = ~n10485 & ~n10486;
  assign n10488 = ~n10480 & ~n10487;
  assign n10489 = ~n8241 & ~n10485;
  assign n10490 = ~n10486 & n10489;
  assign n10491 = ~n10479 & n10490;
  assign n10492 = ~n10488 & ~n10491;
  assign n10493 = n8203 & ~n8209;
  assign n10494 = ~n8213 & ~n10493;
  assign n10495 = ~n7881 & ~n7898;
  assign n10496 = ~n7894 & ~n10495;
  assign n10497 = ~n7917 & ~n7934;
  assign n10498 = ~n7930 & ~n10497;
  assign n10499 = ~n10496 & n10498;
  assign n10500 = n10496 & ~n10498;
  assign n10501 = ~n10499 & ~n10500;
  assign n10502 = ~n10494 & ~n10501;
  assign n10503 = ~n8213 & ~n10499;
  assign n10504 = ~n10500 & n10503;
  assign n10505 = ~n10493 & n10504;
  assign n10506 = ~n10502 & ~n10505;
  assign n10507 = ~n10492 & n10506;
  assign n10508 = n10492 & ~n10506;
  assign n10509 = ~n10507 & ~n10508;
  assign n10510 = ~n10478 & ~n10509;
  assign n10511 = n10478 & n10509;
  assign n10512 = ~n10510 & ~n10511;
  assign n10513 = ~n8165 & ~n8186;
  assign n10514 = ~n8188 & ~n10513;
  assign n10515 = n8148 & ~n8158;
  assign n10516 = ~n8162 & ~n10515;
  assign n10517 = ~n7803 & ~n7820;
  assign n10518 = ~n7816 & ~n10517;
  assign n10519 = ~n7839 & ~n7856;
  assign n10520 = ~n7852 & ~n10519;
  assign n10521 = ~n10518 & n10520;
  assign n10522 = n10518 & ~n10520;
  assign n10523 = ~n10521 & ~n10522;
  assign n10524 = ~n10516 & ~n10523;
  assign n10525 = ~n8162 & ~n10521;
  assign n10526 = ~n10522 & n10525;
  assign n10527 = ~n10515 & n10526;
  assign n10528 = ~n10524 & ~n10527;
  assign n10529 = n8167 & ~n8173;
  assign n10530 = ~n8177 & ~n10529;
  assign n10531 = ~n7728 & ~n7745;
  assign n10532 = ~n7741 & ~n10531;
  assign n10533 = ~n7764 & ~n7781;
  assign n10534 = ~n7777 & ~n10533;
  assign n10535 = ~n10532 & n10534;
  assign n10536 = n10532 & ~n10534;
  assign n10537 = ~n10535 & ~n10536;
  assign n10538 = ~n10530 & ~n10537;
  assign n10539 = ~n8177 & ~n10535;
  assign n10540 = ~n10536 & n10539;
  assign n10541 = ~n10529 & n10540;
  assign n10542 = ~n10538 & ~n10541;
  assign n10543 = ~n10528 & n10542;
  assign n10544 = n10528 & ~n10542;
  assign n10545 = ~n10543 & ~n10544;
  assign n10546 = ~n10514 & ~n10545;
  assign n10547 = n10514 & n10545;
  assign n10548 = ~n10546 & ~n10547;
  assign n10549 = ~n10512 & n10548;
  assign n10550 = n10512 & ~n10548;
  assign n10551 = ~n10549 & ~n10550;
  assign n10552 = ~n10476 & ~n10551;
  assign n10553 = n10476 & n10551;
  assign n10554 = ~n10552 & ~n10553;
  assign n10555 = ~n8079 & ~n8131;
  assign n10556 = ~n8133 & ~n10555;
  assign n10557 = ~n8072 & ~n8075;
  assign n10558 = ~n8076 & ~n10557;
  assign n10559 = n8055 & ~n8065;
  assign n10560 = ~n8069 & ~n10559;
  assign n10561 = ~n7647 & ~n7664;
  assign n10562 = ~n7660 & ~n10561;
  assign n10563 = ~n7683 & ~n7700;
  assign n10564 = ~n7696 & ~n10563;
  assign n10565 = ~n10562 & n10564;
  assign n10566 = n10562 & ~n10564;
  assign n10567 = ~n10565 & ~n10566;
  assign n10568 = ~n10560 & ~n10567;
  assign n10569 = ~n8069 & ~n10565;
  assign n10570 = ~n10566 & n10569;
  assign n10571 = ~n10559 & n10570;
  assign n10572 = ~n10568 & ~n10571;
  assign n10573 = n8031 & ~n8037;
  assign n10574 = ~n8041 & ~n10573;
  assign n10575 = ~n7572 & ~n7589;
  assign n10576 = ~n7585 & ~n10575;
  assign n10577 = ~n7608 & ~n7625;
  assign n10578 = ~n7621 & ~n10577;
  assign n10579 = ~n10576 & n10578;
  assign n10580 = n10576 & ~n10578;
  assign n10581 = ~n10579 & ~n10580;
  assign n10582 = ~n10574 & ~n10581;
  assign n10583 = ~n8041 & ~n10579;
  assign n10584 = ~n10580 & n10583;
  assign n10585 = ~n10573 & n10584;
  assign n10586 = ~n10582 & ~n10585;
  assign n10587 = ~n10572 & n10586;
  assign n10588 = n10572 & ~n10586;
  assign n10589 = ~n10587 & ~n10588;
  assign n10590 = ~n10558 & ~n10589;
  assign n10591 = n10558 & n10589;
  assign n10592 = ~n10590 & ~n10591;
  assign n10593 = ~n8098 & ~n8119;
  assign n10594 = ~n8121 & ~n10593;
  assign n10595 = n8081 & ~n8091;
  assign n10596 = ~n8095 & ~n10595;
  assign n10597 = ~n7494 & ~n7511;
  assign n10598 = ~n7507 & ~n10597;
  assign n10599 = ~n7530 & ~n7547;
  assign n10600 = ~n7543 & ~n10599;
  assign n10601 = ~n10598 & n10600;
  assign n10602 = n10598 & ~n10600;
  assign n10603 = ~n10601 & ~n10602;
  assign n10604 = ~n10596 & ~n10603;
  assign n10605 = ~n8095 & ~n10601;
  assign n10606 = ~n10602 & n10605;
  assign n10607 = ~n10595 & n10606;
  assign n10608 = ~n10604 & ~n10607;
  assign n10609 = n8100 & ~n8106;
  assign n10610 = ~n8110 & ~n10609;
  assign n10611 = ~n7419 & ~n7436;
  assign n10612 = ~n7432 & ~n10611;
  assign n10613 = ~n7455 & ~n7472;
  assign n10614 = ~n7468 & ~n10613;
  assign n10615 = ~n10612 & n10614;
  assign n10616 = n10612 & ~n10614;
  assign n10617 = ~n10615 & ~n10616;
  assign n10618 = ~n10610 & ~n10617;
  assign n10619 = ~n8110 & ~n10615;
  assign n10620 = ~n10616 & n10619;
  assign n10621 = ~n10609 & n10620;
  assign n10622 = ~n10618 & ~n10621;
  assign n10623 = ~n10608 & n10622;
  assign n10624 = n10608 & ~n10622;
  assign n10625 = ~n10623 & ~n10624;
  assign n10626 = ~n10594 & ~n10625;
  assign n10627 = n10594 & n10625;
  assign n10628 = ~n10626 & ~n10627;
  assign n10629 = ~n10592 & n10628;
  assign n10630 = n10592 & ~n10628;
  assign n10631 = ~n10629 & ~n10630;
  assign n10632 = ~n10556 & ~n10631;
  assign n10633 = n10556 & n10631;
  assign n10634 = ~n10632 & ~n10633;
  assign n10635 = ~n10554 & n10634;
  assign n10636 = n10554 & ~n10634;
  assign n10637 = ~n10635 & ~n10636;
  assign n10638 = ~n10474 & ~n10637;
  assign n10639 = n10474 & n10637;
  assign n10640 = ~n10638 & ~n10639;
  assign n10641 = ~n6964 & ~n7390;
  assign n10642 = ~n7392 & ~n10641;
  assign n10643 = ~n6957 & ~n6960;
  assign n10644 = ~n6961 & ~n10643;
  assign n10645 = ~n6950 & ~n6953;
  assign n10646 = ~n6954 & ~n10645;
  assign n10647 = n6933 & ~n6943;
  assign n10648 = ~n6947 & ~n10647;
  assign n10649 = ~n6840 & ~n6857;
  assign n10650 = ~n6853 & ~n10649;
  assign n10651 = ~n6876 & ~n6893;
  assign n10652 = ~n6889 & ~n10651;
  assign n10653 = ~n10650 & n10652;
  assign n10654 = n10650 & ~n10652;
  assign n10655 = ~n10653 & ~n10654;
  assign n10656 = ~n10648 & ~n10655;
  assign n10657 = ~n6947 & ~n10653;
  assign n10658 = ~n10654 & n10657;
  assign n10659 = ~n10647 & n10658;
  assign n10660 = ~n10656 & ~n10659;
  assign n10661 = n6909 & ~n6915;
  assign n10662 = ~n6919 & ~n10661;
  assign n10663 = ~n6765 & ~n6782;
  assign n10664 = ~n6778 & ~n10663;
  assign n10665 = ~n6801 & ~n6818;
  assign n10666 = ~n6814 & ~n10665;
  assign n10667 = ~n10664 & n10666;
  assign n10668 = n10664 & ~n10666;
  assign n10669 = ~n10667 & ~n10668;
  assign n10670 = ~n10662 & ~n10669;
  assign n10671 = ~n6919 & ~n10667;
  assign n10672 = ~n10668 & n10671;
  assign n10673 = ~n10661 & n10672;
  assign n10674 = ~n10670 & ~n10673;
  assign n10675 = ~n10660 & n10674;
  assign n10676 = n10660 & ~n10674;
  assign n10677 = ~n10675 & ~n10676;
  assign n10678 = ~n10646 & ~n10677;
  assign n10679 = n10646 & n10677;
  assign n10680 = ~n10678 & ~n10679;
  assign n10681 = ~n6635 & ~n6736;
  assign n10682 = ~n6738 & ~n10681;
  assign n10683 = n6582 & ~n6628;
  assign n10684 = ~n6632 & ~n10683;
  assign n10685 = ~n6614 & ~n6618;
  assign n10686 = ~n6610 & ~n10685;
  assign n10687 = ~n6574 & ~n6577;
  assign n10688 = ~n6580 & ~n10687;
  assign n10689 = ~n10686 & n10688;
  assign n10690 = n10686 & ~n10688;
  assign n10691 = ~n10689 & ~n10690;
  assign n10692 = ~n10684 & ~n10691;
  assign n10693 = ~n6632 & ~n10689;
  assign n10694 = ~n10690 & n10693;
  assign n10695 = ~n10683 & n10694;
  assign n10696 = ~n10692 & ~n10695;
  assign n10697 = n6671 & ~n6713;
  assign n10698 = ~n6717 & ~n10697;
  assign n10699 = ~n6703 & ~n6707;
  assign n10700 = ~n6699 & ~n10699;
  assign n10701 = ~n6663 & ~n6666;
  assign n10702 = ~n6669 & ~n10701;
  assign n10703 = ~n10700 & n10702;
  assign n10704 = n10700 & ~n10702;
  assign n10705 = ~n10703 & ~n10704;
  assign n10706 = ~n10698 & ~n10705;
  assign n10707 = ~n6717 & ~n10703;
  assign n10708 = ~n10704 & n10707;
  assign n10709 = ~n10697 & n10708;
  assign n10710 = ~n10706 & ~n10709;
  assign n10711 = ~n10696 & n10710;
  assign n10712 = n10696 & ~n10710;
  assign n10713 = ~n10711 & ~n10712;
  assign n10714 = ~n10682 & ~n10713;
  assign n10715 = n10682 & n10713;
  assign n10716 = ~n10714 & ~n10715;
  assign n10717 = ~n10680 & n10716;
  assign n10718 = n10680 & ~n10716;
  assign n10719 = ~n10717 & ~n10718;
  assign n10720 = ~n10644 & ~n10719;
  assign n10721 = n10644 & n10719;
  assign n10722 = ~n10720 & ~n10721;
  assign n10723 = ~n7164 & ~n7372;
  assign n10724 = ~n7374 & ~n10723;
  assign n10725 = ~n7157 & ~n7160;
  assign n10726 = ~n7161 & ~n10725;
  assign n10727 = n7140 & ~n7150;
  assign n10728 = ~n7154 & ~n10727;
  assign n10729 = ~n7074 & ~n7091;
  assign n10730 = ~n7087 & ~n10729;
  assign n10731 = ~n7110 & ~n7127;
  assign n10732 = ~n7123 & ~n10731;
  assign n10733 = ~n10730 & n10732;
  assign n10734 = n10730 & ~n10732;
  assign n10735 = ~n10733 & ~n10734;
  assign n10736 = ~n10728 & ~n10735;
  assign n10737 = ~n7154 & ~n10733;
  assign n10738 = ~n10734 & n10737;
  assign n10739 = ~n10727 & n10738;
  assign n10740 = ~n10736 & ~n10739;
  assign n10741 = n7000 & ~n7042;
  assign n10742 = ~n7046 & ~n10741;
  assign n10743 = ~n7032 & ~n7036;
  assign n10744 = ~n7028 & ~n10743;
  assign n10745 = ~n6992 & ~n6995;
  assign n10746 = ~n6998 & ~n10745;
  assign n10747 = ~n10744 & n10746;
  assign n10748 = n10744 & ~n10746;
  assign n10749 = ~n10747 & ~n10748;
  assign n10750 = ~n10742 & ~n10749;
  assign n10751 = ~n7046 & ~n10747;
  assign n10752 = ~n10748 & n10751;
  assign n10753 = ~n10741 & n10752;
  assign n10754 = ~n10750 & ~n10753;
  assign n10755 = ~n10740 & n10754;
  assign n10756 = n10740 & ~n10754;
  assign n10757 = ~n10755 & ~n10756;
  assign n10758 = ~n10726 & ~n10757;
  assign n10759 = n10726 & n10757;
  assign n10760 = ~n10758 & ~n10759;
  assign n10761 = ~n7253 & ~n7354;
  assign n10762 = ~n7356 & ~n10761;
  assign n10763 = n7200 & ~n7246;
  assign n10764 = ~n7250 & ~n10763;
  assign n10765 = ~n7232 & ~n7236;
  assign n10766 = ~n7228 & ~n10765;
  assign n10767 = ~n7192 & ~n7195;
  assign n10768 = ~n7198 & ~n10767;
  assign n10769 = ~n10766 & n10768;
  assign n10770 = n10766 & ~n10768;
  assign n10771 = ~n10769 & ~n10770;
  assign n10772 = ~n10764 & ~n10771;
  assign n10773 = ~n7250 & ~n10769;
  assign n10774 = ~n10770 & n10773;
  assign n10775 = ~n10763 & n10774;
  assign n10776 = ~n10772 & ~n10775;
  assign n10777 = n7289 & ~n7331;
  assign n10778 = ~n7335 & ~n10777;
  assign n10779 = ~n7321 & ~n7325;
  assign n10780 = ~n7317 & ~n10779;
  assign n10781 = ~n7281 & ~n7284;
  assign n10782 = ~n7287 & ~n10781;
  assign n10783 = ~n10780 & n10782;
  assign n10784 = n10780 & ~n10782;
  assign n10785 = ~n10783 & ~n10784;
  assign n10786 = ~n10778 & ~n10785;
  assign n10787 = ~n7335 & ~n10783;
  assign n10788 = ~n10784 & n10787;
  assign n10789 = ~n10777 & n10788;
  assign n10790 = ~n10786 & ~n10789;
  assign n10791 = ~n10776 & n10790;
  assign n10792 = n10776 & ~n10790;
  assign n10793 = ~n10791 & ~n10792;
  assign n10794 = ~n10762 & ~n10793;
  assign n10795 = n10762 & n10793;
  assign n10796 = ~n10794 & ~n10795;
  assign n10797 = ~n10760 & n10796;
  assign n10798 = n10760 & ~n10796;
  assign n10799 = ~n10797 & ~n10798;
  assign n10800 = ~n10724 & ~n10799;
  assign n10801 = n10724 & n10799;
  assign n10802 = ~n10800 & ~n10801;
  assign n10803 = ~n10722 & n10802;
  assign n10804 = n10722 & ~n10802;
  assign n10805 = ~n10803 & ~n10804;
  assign n10806 = ~n10642 & ~n10805;
  assign n10807 = n10642 & n10805;
  assign n10808 = ~n10806 & ~n10807;
  assign n10809 = ~n10640 & n10808;
  assign n10810 = n10640 & ~n10808;
  assign n10811 = ~n10809 & ~n10810;
  assign n10812 = ~n10472 & ~n10811;
  assign n10813 = n10472 & n10811;
  assign n10814 = ~n10812 & ~n10813;
  assign n10815 = ~n9126 & ~n9988;
  assign n10816 = ~n9990 & ~n10815;
  assign n10817 = ~n9119 & ~n9122;
  assign n10818 = ~n9123 & ~n10817;
  assign n10819 = ~n9112 & ~n9115;
  assign n10820 = ~n9116 & ~n10819;
  assign n10821 = ~n9105 & ~n9108;
  assign n10822 = ~n9109 & ~n10821;
  assign n10823 = n9088 & ~n9098;
  assign n10824 = ~n9102 & ~n10823;
  assign n10825 = ~n8937 & ~n8954;
  assign n10826 = ~n8950 & ~n10825;
  assign n10827 = ~n8973 & ~n8990;
  assign n10828 = ~n8986 & ~n10827;
  assign n10829 = ~n10826 & n10828;
  assign n10830 = n10826 & ~n10828;
  assign n10831 = ~n10829 & ~n10830;
  assign n10832 = ~n10824 & ~n10831;
  assign n10833 = ~n9102 & ~n10829;
  assign n10834 = ~n10830 & n10833;
  assign n10835 = ~n10823 & n10834;
  assign n10836 = ~n10832 & ~n10835;
  assign n10837 = n9064 & ~n9070;
  assign n10838 = ~n9074 & ~n10837;
  assign n10839 = ~n8862 & ~n8879;
  assign n10840 = ~n8875 & ~n10839;
  assign n10841 = ~n8898 & ~n8915;
  assign n10842 = ~n8911 & ~n10841;
  assign n10843 = ~n10840 & n10842;
  assign n10844 = n10840 & ~n10842;
  assign n10845 = ~n10843 & ~n10844;
  assign n10846 = ~n10838 & ~n10845;
  assign n10847 = ~n9074 & ~n10843;
  assign n10848 = ~n10844 & n10847;
  assign n10849 = ~n10837 & n10848;
  assign n10850 = ~n10846 & ~n10849;
  assign n10851 = ~n10836 & n10850;
  assign n10852 = n10836 & ~n10850;
  assign n10853 = ~n10851 & ~n10852;
  assign n10854 = ~n10822 & ~n10853;
  assign n10855 = n10822 & n10853;
  assign n10856 = ~n10854 & ~n10855;
  assign n10857 = ~n9026 & ~n9047;
  assign n10858 = ~n9049 & ~n10857;
  assign n10859 = n9009 & ~n9019;
  assign n10860 = ~n9023 & ~n10859;
  assign n10861 = ~n8784 & ~n8801;
  assign n10862 = ~n8797 & ~n10861;
  assign n10863 = ~n8820 & ~n8837;
  assign n10864 = ~n8833 & ~n10863;
  assign n10865 = ~n10862 & n10864;
  assign n10866 = n10862 & ~n10864;
  assign n10867 = ~n10865 & ~n10866;
  assign n10868 = ~n10860 & ~n10867;
  assign n10869 = ~n9023 & ~n10865;
  assign n10870 = ~n10866 & n10869;
  assign n10871 = ~n10859 & n10870;
  assign n10872 = ~n10868 & ~n10871;
  assign n10873 = n9028 & ~n9034;
  assign n10874 = ~n9038 & ~n10873;
  assign n10875 = ~n8709 & ~n8726;
  assign n10876 = ~n8722 & ~n10875;
  assign n10877 = ~n8745 & ~n8762;
  assign n10878 = ~n8758 & ~n10877;
  assign n10879 = ~n10876 & n10878;
  assign n10880 = n10876 & ~n10878;
  assign n10881 = ~n10879 & ~n10880;
  assign n10882 = ~n10874 & ~n10881;
  assign n10883 = ~n9038 & ~n10879;
  assign n10884 = ~n10880 & n10883;
  assign n10885 = ~n10873 & n10884;
  assign n10886 = ~n10882 & ~n10885;
  assign n10887 = ~n10872 & n10886;
  assign n10888 = n10872 & ~n10886;
  assign n10889 = ~n10887 & ~n10888;
  assign n10890 = ~n10858 & ~n10889;
  assign n10891 = n10858 & n10889;
  assign n10892 = ~n10890 & ~n10891;
  assign n10893 = ~n10856 & n10892;
  assign n10894 = n10856 & ~n10892;
  assign n10895 = ~n10893 & ~n10894;
  assign n10896 = ~n10820 & ~n10895;
  assign n10897 = n10820 & n10895;
  assign n10898 = ~n10896 & ~n10897;
  assign n10899 = ~n8472 & ~n8680;
  assign n10900 = ~n8682 & ~n10899;
  assign n10901 = ~n8465 & ~n8468;
  assign n10902 = ~n8469 & ~n10901;
  assign n10903 = n8448 & ~n8458;
  assign n10904 = ~n8462 & ~n10903;
  assign n10905 = ~n8382 & ~n8399;
  assign n10906 = ~n8395 & ~n10905;
  assign n10907 = ~n8418 & ~n8435;
  assign n10908 = ~n8431 & ~n10907;
  assign n10909 = ~n10906 & n10908;
  assign n10910 = n10906 & ~n10908;
  assign n10911 = ~n10909 & ~n10910;
  assign n10912 = ~n10904 & ~n10911;
  assign n10913 = ~n8462 & ~n10909;
  assign n10914 = ~n10910 & n10913;
  assign n10915 = ~n10903 & n10914;
  assign n10916 = ~n10912 & ~n10915;
  assign n10917 = n8308 & ~n8350;
  assign n10918 = ~n8354 & ~n10917;
  assign n10919 = ~n8340 & ~n8344;
  assign n10920 = ~n8336 & ~n10919;
  assign n10921 = ~n8300 & ~n8303;
  assign n10922 = ~n8306 & ~n10921;
  assign n10923 = ~n10920 & n10922;
  assign n10924 = n10920 & ~n10922;
  assign n10925 = ~n10923 & ~n10924;
  assign n10926 = ~n10918 & ~n10925;
  assign n10927 = ~n8354 & ~n10923;
  assign n10928 = ~n10924 & n10927;
  assign n10929 = ~n10917 & n10928;
  assign n10930 = ~n10926 & ~n10929;
  assign n10931 = ~n10916 & n10930;
  assign n10932 = n10916 & ~n10930;
  assign n10933 = ~n10931 & ~n10932;
  assign n10934 = ~n10902 & ~n10933;
  assign n10935 = n10902 & n10933;
  assign n10936 = ~n10934 & ~n10935;
  assign n10937 = ~n8561 & ~n8662;
  assign n10938 = ~n8664 & ~n10937;
  assign n10939 = n8508 & ~n8554;
  assign n10940 = ~n8558 & ~n10939;
  assign n10941 = ~n8540 & ~n8544;
  assign n10942 = ~n8536 & ~n10941;
  assign n10943 = ~n8500 & ~n8503;
  assign n10944 = ~n8506 & ~n10943;
  assign n10945 = ~n10942 & n10944;
  assign n10946 = n10942 & ~n10944;
  assign n10947 = ~n10945 & ~n10946;
  assign n10948 = ~n10940 & ~n10947;
  assign n10949 = ~n8558 & ~n10945;
  assign n10950 = ~n10946 & n10949;
  assign n10951 = ~n10939 & n10950;
  assign n10952 = ~n10948 & ~n10951;
  assign n10953 = n8597 & ~n8639;
  assign n10954 = ~n8643 & ~n10953;
  assign n10955 = ~n8629 & ~n8633;
  assign n10956 = ~n8625 & ~n10955;
  assign n10957 = ~n8589 & ~n8592;
  assign n10958 = ~n8595 & ~n10957;
  assign n10959 = ~n10956 & n10958;
  assign n10960 = n10956 & ~n10958;
  assign n10961 = ~n10959 & ~n10960;
  assign n10962 = ~n10954 & ~n10961;
  assign n10963 = ~n8643 & ~n10959;
  assign n10964 = ~n10960 & n10963;
  assign n10965 = ~n10953 & n10964;
  assign n10966 = ~n10962 & ~n10965;
  assign n10967 = ~n10952 & n10966;
  assign n10968 = n10952 & ~n10966;
  assign n10969 = ~n10967 & ~n10968;
  assign n10970 = ~n10938 & ~n10969;
  assign n10971 = n10938 & n10969;
  assign n10972 = ~n10970 & ~n10971;
  assign n10973 = ~n10936 & n10972;
  assign n10974 = n10936 & ~n10972;
  assign n10975 = ~n10973 & ~n10974;
  assign n10976 = ~n10900 & ~n10975;
  assign n10977 = n10900 & n10975;
  assign n10978 = ~n10976 & ~n10977;
  assign n10979 = ~n10898 & n10978;
  assign n10980 = n10898 & ~n10978;
  assign n10981 = ~n10979 & ~n10980;
  assign n10982 = ~n10818 & ~n10981;
  assign n10983 = n10818 & n10981;
  assign n10984 = ~n10982 & ~n10983;
  assign n10985 = ~n9544 & ~n9970;
  assign n10986 = ~n9972 & ~n10985;
  assign n10987 = ~n9537 & ~n9540;
  assign n10988 = ~n9541 & ~n10987;
  assign n10989 = ~n9530 & ~n9533;
  assign n10990 = ~n9534 & ~n10989;
  assign n10991 = n9513 & ~n9523;
  assign n10992 = ~n9527 & ~n10991;
  assign n10993 = ~n9420 & ~n9437;
  assign n10994 = ~n9433 & ~n10993;
  assign n10995 = ~n9456 & ~n9473;
  assign n10996 = ~n9469 & ~n10995;
  assign n10997 = ~n10994 & n10996;
  assign n10998 = n10994 & ~n10996;
  assign n10999 = ~n10997 & ~n10998;
  assign n11000 = ~n10992 & ~n10999;
  assign n11001 = ~n9527 & ~n10997;
  assign n11002 = ~n10998 & n11001;
  assign n11003 = ~n10991 & n11002;
  assign n11004 = ~n11000 & ~n11003;
  assign n11005 = n9489 & ~n9495;
  assign n11006 = ~n9499 & ~n11005;
  assign n11007 = ~n9345 & ~n9362;
  assign n11008 = ~n9358 & ~n11007;
  assign n11009 = ~n9381 & ~n9398;
  assign n11010 = ~n9394 & ~n11009;
  assign n11011 = ~n11008 & n11010;
  assign n11012 = n11008 & ~n11010;
  assign n11013 = ~n11011 & ~n11012;
  assign n11014 = ~n11006 & ~n11013;
  assign n11015 = ~n9499 & ~n11011;
  assign n11016 = ~n11012 & n11015;
  assign n11017 = ~n11005 & n11016;
  assign n11018 = ~n11014 & ~n11017;
  assign n11019 = ~n11004 & n11018;
  assign n11020 = n11004 & ~n11018;
  assign n11021 = ~n11019 & ~n11020;
  assign n11022 = ~n10990 & ~n11021;
  assign n11023 = n10990 & n11021;
  assign n11024 = ~n11022 & ~n11023;
  assign n11025 = ~n9215 & ~n9316;
  assign n11026 = ~n9318 & ~n11025;
  assign n11027 = n9162 & ~n9208;
  assign n11028 = ~n9212 & ~n11027;
  assign n11029 = ~n9194 & ~n9198;
  assign n11030 = ~n9190 & ~n11029;
  assign n11031 = ~n9154 & ~n9157;
  assign n11032 = ~n9160 & ~n11031;
  assign n11033 = ~n11030 & n11032;
  assign n11034 = n11030 & ~n11032;
  assign n11035 = ~n11033 & ~n11034;
  assign n11036 = ~n11028 & ~n11035;
  assign n11037 = ~n9212 & ~n11033;
  assign n11038 = ~n11034 & n11037;
  assign n11039 = ~n11027 & n11038;
  assign n11040 = ~n11036 & ~n11039;
  assign n11041 = n9251 & ~n9293;
  assign n11042 = ~n9297 & ~n11041;
  assign n11043 = ~n9283 & ~n9287;
  assign n11044 = ~n9279 & ~n11043;
  assign n11045 = ~n9243 & ~n9246;
  assign n11046 = ~n9249 & ~n11045;
  assign n11047 = ~n11044 & n11046;
  assign n11048 = n11044 & ~n11046;
  assign n11049 = ~n11047 & ~n11048;
  assign n11050 = ~n11042 & ~n11049;
  assign n11051 = ~n9297 & ~n11047;
  assign n11052 = ~n11048 & n11051;
  assign n11053 = ~n11041 & n11052;
  assign n11054 = ~n11050 & ~n11053;
  assign n11055 = ~n11040 & n11054;
  assign n11056 = n11040 & ~n11054;
  assign n11057 = ~n11055 & ~n11056;
  assign n11058 = ~n11026 & ~n11057;
  assign n11059 = n11026 & n11057;
  assign n11060 = ~n11058 & ~n11059;
  assign n11061 = ~n11024 & n11060;
  assign n11062 = n11024 & ~n11060;
  assign n11063 = ~n11061 & ~n11062;
  assign n11064 = ~n10988 & ~n11063;
  assign n11065 = n10988 & n11063;
  assign n11066 = ~n11064 & ~n11065;
  assign n11067 = ~n9744 & ~n9952;
  assign n11068 = ~n9954 & ~n11067;
  assign n11069 = ~n9737 & ~n9740;
  assign n11070 = ~n9741 & ~n11069;
  assign n11071 = n9720 & ~n9730;
  assign n11072 = ~n9734 & ~n11071;
  assign n11073 = ~n9654 & ~n9671;
  assign n11074 = ~n9667 & ~n11073;
  assign n11075 = ~n9690 & ~n9707;
  assign n11076 = ~n9703 & ~n11075;
  assign n11077 = ~n11074 & n11076;
  assign n11078 = n11074 & ~n11076;
  assign n11079 = ~n11077 & ~n11078;
  assign n11080 = ~n11072 & ~n11079;
  assign n11081 = ~n9734 & ~n11077;
  assign n11082 = ~n11078 & n11081;
  assign n11083 = ~n11071 & n11082;
  assign n11084 = ~n11080 & ~n11083;
  assign n11085 = n9580 & ~n9622;
  assign n11086 = ~n9626 & ~n11085;
  assign n11087 = ~n9612 & ~n9616;
  assign n11088 = ~n9608 & ~n11087;
  assign n11089 = ~n9572 & ~n9575;
  assign n11090 = ~n9578 & ~n11089;
  assign n11091 = ~n11088 & n11090;
  assign n11092 = n11088 & ~n11090;
  assign n11093 = ~n11091 & ~n11092;
  assign n11094 = ~n11086 & ~n11093;
  assign n11095 = ~n9626 & ~n11091;
  assign n11096 = ~n11092 & n11095;
  assign n11097 = ~n11085 & n11096;
  assign n11098 = ~n11094 & ~n11097;
  assign n11099 = ~n11084 & n11098;
  assign n11100 = n11084 & ~n11098;
  assign n11101 = ~n11099 & ~n11100;
  assign n11102 = ~n11070 & ~n11101;
  assign n11103 = n11070 & n11101;
  assign n11104 = ~n11102 & ~n11103;
  assign n11105 = ~n9833 & ~n9934;
  assign n11106 = ~n9936 & ~n11105;
  assign n11107 = n9780 & ~n9826;
  assign n11108 = ~n9830 & ~n11107;
  assign n11109 = ~n9812 & ~n9816;
  assign n11110 = ~n9808 & ~n11109;
  assign n11111 = ~n9772 & ~n9775;
  assign n11112 = ~n9778 & ~n11111;
  assign n11113 = ~n11110 & n11112;
  assign n11114 = n11110 & ~n11112;
  assign n11115 = ~n11113 & ~n11114;
  assign n11116 = ~n11108 & ~n11115;
  assign n11117 = ~n9830 & ~n11113;
  assign n11118 = ~n11114 & n11117;
  assign n11119 = ~n11107 & n11118;
  assign n11120 = ~n11116 & ~n11119;
  assign n11121 = n9869 & ~n9911;
  assign n11122 = ~n9915 & ~n11121;
  assign n11123 = ~n9901 & ~n9905;
  assign n11124 = ~n9897 & ~n11123;
  assign n11125 = ~n9861 & ~n9864;
  assign n11126 = ~n9867 & ~n11125;
  assign n11127 = ~n11124 & n11126;
  assign n11128 = n11124 & ~n11126;
  assign n11129 = ~n11127 & ~n11128;
  assign n11130 = ~n11122 & ~n11129;
  assign n11131 = ~n9915 & ~n11127;
  assign n11132 = ~n11128 & n11131;
  assign n11133 = ~n11121 & n11132;
  assign n11134 = ~n11130 & ~n11133;
  assign n11135 = ~n11120 & n11134;
  assign n11136 = n11120 & ~n11134;
  assign n11137 = ~n11135 & ~n11136;
  assign n11138 = ~n11106 & ~n11137;
  assign n11139 = n11106 & n11137;
  assign n11140 = ~n11138 & ~n11139;
  assign n11141 = ~n11104 & n11140;
  assign n11142 = n11104 & ~n11140;
  assign n11143 = ~n11141 & ~n11142;
  assign n11144 = ~n11068 & ~n11143;
  assign n11145 = n11068 & n11143;
  assign n11146 = ~n11144 & ~n11145;
  assign n11147 = ~n11066 & n11146;
  assign n11148 = n11066 & ~n11146;
  assign n11149 = ~n11147 & ~n11148;
  assign n11150 = ~n10986 & ~n11149;
  assign n11151 = n10986 & n11149;
  assign n11152 = ~n11150 & ~n11151;
  assign n11153 = ~n10984 & n11152;
  assign n11154 = n10984 & ~n11152;
  assign n11155 = ~n11153 & ~n11154;
  assign n11156 = ~n10816 & ~n11155;
  assign n11157 = n10816 & n11155;
  assign n11158 = ~n11156 & ~n11157;
  assign n11159 = ~n10814 & n11158;
  assign n11160 = n10814 & ~n11158;
  assign n11161 = ~n11159 & ~n11160;
  assign n11162 = ~n10470 & ~n11161;
  assign n11163 = n10470 & n11161;
  assign n11164 = ~n11162 & ~n11163;
  assign n11165 = ~n10468 & n11164;
  assign n11166 = n10468 & ~n11164;
  assign n11167 = ~n11165 & ~n11166;
  assign n11168 = ~n10049 & ~n11167;
  assign n11169 = n10049 & n11167;
  assign n11170 = ~n11168 & ~n11169;
  assign n11171 = ~n4465 & ~n4468;
  assign n11172 = ~n4469 & ~n11171;
  assign n11173 = ~n4458 & ~n4461;
  assign n11174 = ~n4462 & ~n11173;
  assign n11175 = ~n4451 & ~n4454;
  assign n11176 = ~n4455 & ~n11175;
  assign n11177 = ~n4444 & ~n4447;
  assign n11178 = ~n4448 & ~n11177;
  assign n11179 = ~n4437 & ~n4440;
  assign n11180 = ~n4441 & ~n11179;
  assign n11181 = n4420 & ~n4430;
  assign n11182 = ~n4434 & ~n11181;
  assign n11183 = ~n2744 & ~n2761;
  assign n11184 = ~n2757 & ~n11183;
  assign n11185 = ~n2780 & ~n2794;
  assign n11186 = ~n2797 & ~n11185;
  assign n11187 = ~n11184 & n11186;
  assign n11188 = n11184 & ~n11186;
  assign n11189 = ~n11187 & ~n11188;
  assign n11190 = ~n11182 & ~n11189;
  assign n11191 = ~n4434 & ~n11187;
  assign n11192 = ~n11188 & n11191;
  assign n11193 = ~n11181 & n11192;
  assign n11194 = ~n11190 & ~n11193;
  assign n11195 = n4396 & ~n4402;
  assign n11196 = ~n4406 & ~n11195;
  assign n11197 = ~n2819 & ~n2836;
  assign n11198 = ~n2832 & ~n11197;
  assign n11199 = ~n2855 & ~n2872;
  assign n11200 = ~n2868 & ~n11199;
  assign n11201 = ~n11198 & n11200;
  assign n11202 = n11198 & ~n11200;
  assign n11203 = ~n11201 & ~n11202;
  assign n11204 = ~n11196 & ~n11203;
  assign n11205 = ~n4406 & ~n11201;
  assign n11206 = ~n11202 & n11205;
  assign n11207 = ~n11195 & n11206;
  assign n11208 = ~n11204 & ~n11207;
  assign n11209 = ~n11194 & n11208;
  assign n11210 = n11194 & ~n11208;
  assign n11211 = ~n11209 & ~n11210;
  assign n11212 = ~n11180 & ~n11211;
  assign n11213 = n11180 & n11211;
  assign n11214 = ~n11212 & ~n11213;
  assign n11215 = ~n4358 & ~n4379;
  assign n11216 = ~n4381 & ~n11215;
  assign n11217 = n4341 & ~n4351;
  assign n11218 = ~n4355 & ~n11217;
  assign n11219 = ~n2972 & ~n2989;
  assign n11220 = ~n2985 & ~n11219;
  assign n11221 = ~n3008 & ~n3025;
  assign n11222 = ~n3021 & ~n11221;
  assign n11223 = ~n11220 & n11222;
  assign n11224 = n11220 & ~n11222;
  assign n11225 = ~n11223 & ~n11224;
  assign n11226 = ~n11218 & ~n11225;
  assign n11227 = ~n4355 & ~n11223;
  assign n11228 = ~n11224 & n11227;
  assign n11229 = ~n11217 & n11228;
  assign n11230 = ~n11226 & ~n11229;
  assign n11231 = n4360 & ~n4366;
  assign n11232 = ~n4370 & ~n11231;
  assign n11233 = ~n2897 & ~n2914;
  assign n11234 = ~n2910 & ~n11233;
  assign n11235 = ~n2933 & ~n2950;
  assign n11236 = ~n2946 & ~n11235;
  assign n11237 = ~n11234 & n11236;
  assign n11238 = n11234 & ~n11236;
  assign n11239 = ~n11237 & ~n11238;
  assign n11240 = ~n11232 & ~n11239;
  assign n11241 = ~n4370 & ~n11237;
  assign n11242 = ~n11238 & n11241;
  assign n11243 = ~n11231 & n11242;
  assign n11244 = ~n11240 & ~n11243;
  assign n11245 = ~n11230 & n11244;
  assign n11246 = n11230 & ~n11244;
  assign n11247 = ~n11245 & ~n11246;
  assign n11248 = ~n11216 & ~n11247;
  assign n11249 = n11216 & n11247;
  assign n11250 = ~n11248 & ~n11249;
  assign n11251 = ~n11214 & n11250;
  assign n11252 = n11214 & ~n11250;
  assign n11253 = ~n11251 & ~n11252;
  assign n11254 = ~n11178 & ~n11253;
  assign n11255 = n11178 & n11253;
  assign n11256 = ~n11254 & ~n11255;
  assign n11257 = ~n4272 & ~n4324;
  assign n11258 = ~n4326 & ~n11257;
  assign n11259 = ~n4265 & ~n4268;
  assign n11260 = ~n4269 & ~n11259;
  assign n11261 = n4248 & ~n4258;
  assign n11262 = ~n4262 & ~n11261;
  assign n11263 = ~n3281 & ~n3298;
  assign n11264 = ~n3294 & ~n11263;
  assign n11265 = ~n3317 & ~n3334;
  assign n11266 = ~n3330 & ~n11265;
  assign n11267 = ~n11264 & n11266;
  assign n11268 = n11264 & ~n11266;
  assign n11269 = ~n11267 & ~n11268;
  assign n11270 = ~n11262 & ~n11269;
  assign n11271 = ~n4262 & ~n11267;
  assign n11272 = ~n11268 & n11271;
  assign n11273 = ~n11261 & n11272;
  assign n11274 = ~n11270 & ~n11273;
  assign n11275 = n4224 & ~n4230;
  assign n11276 = ~n4234 & ~n11275;
  assign n11277 = ~n3206 & ~n3223;
  assign n11278 = ~n3219 & ~n11277;
  assign n11279 = ~n3242 & ~n3259;
  assign n11280 = ~n3255 & ~n11279;
  assign n11281 = ~n11278 & n11280;
  assign n11282 = n11278 & ~n11280;
  assign n11283 = ~n11281 & ~n11282;
  assign n11284 = ~n11276 & ~n11283;
  assign n11285 = ~n4234 & ~n11281;
  assign n11286 = ~n11282 & n11285;
  assign n11287 = ~n11275 & n11286;
  assign n11288 = ~n11284 & ~n11287;
  assign n11289 = ~n11274 & n11288;
  assign n11290 = n11274 & ~n11288;
  assign n11291 = ~n11289 & ~n11290;
  assign n11292 = ~n11260 & ~n11291;
  assign n11293 = n11260 & n11291;
  assign n11294 = ~n11292 & ~n11293;
  assign n11295 = ~n4291 & ~n4312;
  assign n11296 = ~n4314 & ~n11295;
  assign n11297 = n4274 & ~n4284;
  assign n11298 = ~n4288 & ~n11297;
  assign n11299 = ~n3128 & ~n3145;
  assign n11300 = ~n3141 & ~n11299;
  assign n11301 = ~n3164 & ~n3181;
  assign n11302 = ~n3177 & ~n11301;
  assign n11303 = ~n11300 & n11302;
  assign n11304 = n11300 & ~n11302;
  assign n11305 = ~n11303 & ~n11304;
  assign n11306 = ~n11298 & ~n11305;
  assign n11307 = ~n4288 & ~n11303;
  assign n11308 = ~n11304 & n11307;
  assign n11309 = ~n11297 & n11308;
  assign n11310 = ~n11306 & ~n11309;
  assign n11311 = n4293 & ~n4299;
  assign n11312 = ~n4303 & ~n11311;
  assign n11313 = ~n3053 & ~n3070;
  assign n11314 = ~n3066 & ~n11313;
  assign n11315 = ~n3089 & ~n3106;
  assign n11316 = ~n3102 & ~n11315;
  assign n11317 = ~n11314 & n11316;
  assign n11318 = n11314 & ~n11316;
  assign n11319 = ~n11317 & ~n11318;
  assign n11320 = ~n11312 & ~n11319;
  assign n11321 = ~n4303 & ~n11317;
  assign n11322 = ~n11318 & n11321;
  assign n11323 = ~n11311 & n11322;
  assign n11324 = ~n11320 & ~n11323;
  assign n11325 = ~n11310 & n11324;
  assign n11326 = n11310 & ~n11324;
  assign n11327 = ~n11325 & ~n11326;
  assign n11328 = ~n11296 & ~n11327;
  assign n11329 = n11296 & n11327;
  assign n11330 = ~n11328 & ~n11329;
  assign n11331 = ~n11294 & n11330;
  assign n11332 = n11294 & ~n11330;
  assign n11333 = ~n11331 & ~n11332;
  assign n11334 = ~n11258 & ~n11333;
  assign n11335 = n11258 & n11333;
  assign n11336 = ~n11334 & ~n11335;
  assign n11337 = ~n11256 & n11336;
  assign n11338 = n11256 & ~n11336;
  assign n11339 = ~n11337 & ~n11338;
  assign n11340 = ~n11176 & ~n11339;
  assign n11341 = n11176 & n11339;
  assign n11342 = ~n11340 & ~n11341;
  assign n11343 = ~n4093 & ~n4207;
  assign n11344 = ~n4209 & ~n11343;
  assign n11345 = ~n4086 & ~n4089;
  assign n11346 = ~n4090 & ~n11345;
  assign n11347 = ~n4079 & ~n4082;
  assign n11348 = ~n4083 & ~n11347;
  assign n11349 = n4062 & ~n4072;
  assign n11350 = ~n4076 & ~n11349;
  assign n11351 = ~n3902 & ~n3919;
  assign n11352 = ~n3915 & ~n11351;
  assign n11353 = ~n3938 & ~n3955;
  assign n11354 = ~n3951 & ~n11353;
  assign n11355 = ~n11352 & n11354;
  assign n11356 = n11352 & ~n11354;
  assign n11357 = ~n11355 & ~n11356;
  assign n11358 = ~n11350 & ~n11357;
  assign n11359 = ~n4076 & ~n11355;
  assign n11360 = ~n11356 & n11359;
  assign n11361 = ~n11349 & n11360;
  assign n11362 = ~n11358 & ~n11361;
  assign n11363 = n4038 & ~n4044;
  assign n11364 = ~n4048 & ~n11363;
  assign n11365 = ~n3827 & ~n3844;
  assign n11366 = ~n3840 & ~n11365;
  assign n11367 = ~n3863 & ~n3880;
  assign n11368 = ~n3876 & ~n11367;
  assign n11369 = ~n11366 & n11368;
  assign n11370 = n11366 & ~n11368;
  assign n11371 = ~n11369 & ~n11370;
  assign n11372 = ~n11364 & ~n11371;
  assign n11373 = ~n4048 & ~n11369;
  assign n11374 = ~n11370 & n11373;
  assign n11375 = ~n11363 & n11374;
  assign n11376 = ~n11372 & ~n11375;
  assign n11377 = ~n11362 & n11376;
  assign n11378 = n11362 & ~n11376;
  assign n11379 = ~n11377 & ~n11378;
  assign n11380 = ~n11348 & ~n11379;
  assign n11381 = n11348 & n11379;
  assign n11382 = ~n11380 & ~n11381;
  assign n11383 = ~n4000 & ~n4021;
  assign n11384 = ~n4023 & ~n11383;
  assign n11385 = n3983 & ~n3993;
  assign n11386 = ~n3997 & ~n11385;
  assign n11387 = ~n3749 & ~n3766;
  assign n11388 = ~n3762 & ~n11387;
  assign n11389 = ~n3785 & ~n3802;
  assign n11390 = ~n3798 & ~n11389;
  assign n11391 = ~n11388 & n11390;
  assign n11392 = n11388 & ~n11390;
  assign n11393 = ~n11391 & ~n11392;
  assign n11394 = ~n11386 & ~n11393;
  assign n11395 = ~n3997 & ~n11391;
  assign n11396 = ~n11392 & n11395;
  assign n11397 = ~n11385 & n11396;
  assign n11398 = ~n11394 & ~n11397;
  assign n11399 = n4002 & ~n4008;
  assign n11400 = ~n4012 & ~n11399;
  assign n11401 = ~n3674 & ~n3691;
  assign n11402 = ~n3687 & ~n11401;
  assign n11403 = ~n3710 & ~n3727;
  assign n11404 = ~n3723 & ~n11403;
  assign n11405 = ~n11402 & n11404;
  assign n11406 = n11402 & ~n11404;
  assign n11407 = ~n11405 & ~n11406;
  assign n11408 = ~n11400 & ~n11407;
  assign n11409 = ~n4012 & ~n11405;
  assign n11410 = ~n11406 & n11409;
  assign n11411 = ~n11399 & n11410;
  assign n11412 = ~n11408 & ~n11411;
  assign n11413 = ~n11398 & n11412;
  assign n11414 = n11398 & ~n11412;
  assign n11415 = ~n11413 & ~n11414;
  assign n11416 = ~n11384 & ~n11415;
  assign n11417 = n11384 & n11415;
  assign n11418 = ~n11416 & ~n11417;
  assign n11419 = ~n11382 & n11418;
  assign n11420 = n11382 & ~n11418;
  assign n11421 = ~n11419 & ~n11420;
  assign n11422 = ~n11346 & ~n11421;
  assign n11423 = n11346 & n11421;
  assign n11424 = ~n11422 & ~n11423;
  assign n11425 = ~n4143 & ~n4195;
  assign n11426 = ~n4197 & ~n11425;
  assign n11427 = ~n4136 & ~n4139;
  assign n11428 = ~n4140 & ~n11427;
  assign n11429 = n4119 & ~n4129;
  assign n11430 = ~n4133 & ~n11429;
  assign n11431 = ~n3593 & ~n3610;
  assign n11432 = ~n3606 & ~n11431;
  assign n11433 = ~n3629 & ~n3646;
  assign n11434 = ~n3642 & ~n11433;
  assign n11435 = ~n11432 & n11434;
  assign n11436 = n11432 & ~n11434;
  assign n11437 = ~n11435 & ~n11436;
  assign n11438 = ~n11430 & ~n11437;
  assign n11439 = ~n4133 & ~n11435;
  assign n11440 = ~n11436 & n11439;
  assign n11441 = ~n11429 & n11440;
  assign n11442 = ~n11438 & ~n11441;
  assign n11443 = n4095 & ~n4101;
  assign n11444 = ~n4105 & ~n11443;
  assign n11445 = ~n3518 & ~n3535;
  assign n11446 = ~n3531 & ~n11445;
  assign n11447 = ~n3554 & ~n3571;
  assign n11448 = ~n3567 & ~n11447;
  assign n11449 = ~n11446 & n11448;
  assign n11450 = n11446 & ~n11448;
  assign n11451 = ~n11449 & ~n11450;
  assign n11452 = ~n11444 & ~n11451;
  assign n11453 = ~n4105 & ~n11449;
  assign n11454 = ~n11450 & n11453;
  assign n11455 = ~n11443 & n11454;
  assign n11456 = ~n11452 & ~n11455;
  assign n11457 = ~n11442 & n11456;
  assign n11458 = n11442 & ~n11456;
  assign n11459 = ~n11457 & ~n11458;
  assign n11460 = ~n11428 & ~n11459;
  assign n11461 = n11428 & n11459;
  assign n11462 = ~n11460 & ~n11461;
  assign n11463 = ~n4162 & ~n4183;
  assign n11464 = ~n4185 & ~n11463;
  assign n11465 = n4145 & ~n4155;
  assign n11466 = ~n4159 & ~n11465;
  assign n11467 = ~n3440 & ~n3457;
  assign n11468 = ~n3453 & ~n11467;
  assign n11469 = ~n3476 & ~n3493;
  assign n11470 = ~n3489 & ~n11469;
  assign n11471 = ~n11468 & n11470;
  assign n11472 = n11468 & ~n11470;
  assign n11473 = ~n11471 & ~n11472;
  assign n11474 = ~n11466 & ~n11473;
  assign n11475 = ~n4159 & ~n11471;
  assign n11476 = ~n11472 & n11475;
  assign n11477 = ~n11465 & n11476;
  assign n11478 = ~n11474 & ~n11477;
  assign n11479 = n4164 & ~n4170;
  assign n11480 = ~n4174 & ~n11479;
  assign n11481 = ~n3365 & ~n3382;
  assign n11482 = ~n3378 & ~n11481;
  assign n11483 = ~n3401 & ~n3418;
  assign n11484 = ~n3414 & ~n11483;
  assign n11485 = ~n11482 & n11484;
  assign n11486 = n11482 & ~n11484;
  assign n11487 = ~n11485 & ~n11486;
  assign n11488 = ~n11480 & ~n11487;
  assign n11489 = ~n4174 & ~n11485;
  assign n11490 = ~n11486 & n11489;
  assign n11491 = ~n11479 & n11490;
  assign n11492 = ~n11488 & ~n11491;
  assign n11493 = ~n11478 & n11492;
  assign n11494 = n11478 & ~n11492;
  assign n11495 = ~n11493 & ~n11494;
  assign n11496 = ~n11464 & ~n11495;
  assign n11497 = n11464 & n11495;
  assign n11498 = ~n11496 & ~n11497;
  assign n11499 = ~n11462 & n11498;
  assign n11500 = n11462 & ~n11498;
  assign n11501 = ~n11499 & ~n11500;
  assign n11502 = ~n11426 & ~n11501;
  assign n11503 = n11426 & n11501;
  assign n11504 = ~n11502 & ~n11503;
  assign n11505 = ~n11424 & n11504;
  assign n11506 = n11424 & ~n11504;
  assign n11507 = ~n11505 & ~n11506;
  assign n11508 = ~n11344 & ~n11507;
  assign n11509 = n11344 & n11507;
  assign n11510 = ~n11508 & ~n11509;
  assign n11511 = ~n11342 & n11510;
  assign n11512 = n11342 & ~n11510;
  assign n11513 = ~n11511 & ~n11512;
  assign n11514 = ~n11174 & ~n11513;
  assign n11515 = n11174 & n11513;
  assign n11516 = ~n11514 & ~n11515;
  assign n11517 = ~n1856 & ~n2718;
  assign n11518 = ~n2720 & ~n11517;
  assign n11519 = ~n1849 & ~n1852;
  assign n11520 = ~n1853 & ~n11519;
  assign n11521 = ~n1842 & ~n1845;
  assign n11522 = ~n1846 & ~n11521;
  assign n11523 = ~n1835 & ~n1838;
  assign n11524 = ~n1839 & ~n11523;
  assign n11525 = n1818 & ~n1828;
  assign n11526 = ~n1832 & ~n11525;
  assign n11527 = ~n1667 & ~n1684;
  assign n11528 = ~n1680 & ~n11527;
  assign n11529 = ~n1703 & ~n1720;
  assign n11530 = ~n1716 & ~n11529;
  assign n11531 = ~n11528 & n11530;
  assign n11532 = n11528 & ~n11530;
  assign n11533 = ~n11531 & ~n11532;
  assign n11534 = ~n11526 & ~n11533;
  assign n11535 = ~n1832 & ~n11531;
  assign n11536 = ~n11532 & n11535;
  assign n11537 = ~n11525 & n11536;
  assign n11538 = ~n11534 & ~n11537;
  assign n11539 = n1794 & ~n1800;
  assign n11540 = ~n1804 & ~n11539;
  assign n11541 = ~n1592 & ~n1609;
  assign n11542 = ~n1605 & ~n11541;
  assign n11543 = ~n1628 & ~n1645;
  assign n11544 = ~n1641 & ~n11543;
  assign n11545 = ~n11542 & n11544;
  assign n11546 = n11542 & ~n11544;
  assign n11547 = ~n11545 & ~n11546;
  assign n11548 = ~n11540 & ~n11547;
  assign n11549 = ~n1804 & ~n11545;
  assign n11550 = ~n11546 & n11549;
  assign n11551 = ~n11539 & n11550;
  assign n11552 = ~n11548 & ~n11551;
  assign n11553 = ~n11538 & n11552;
  assign n11554 = n11538 & ~n11552;
  assign n11555 = ~n11553 & ~n11554;
  assign n11556 = ~n11524 & ~n11555;
  assign n11557 = n11524 & n11555;
  assign n11558 = ~n11556 & ~n11557;
  assign n11559 = ~n1756 & ~n1777;
  assign n11560 = ~n1779 & ~n11559;
  assign n11561 = n1739 & ~n1749;
  assign n11562 = ~n1753 & ~n11561;
  assign n11563 = ~n1514 & ~n1531;
  assign n11564 = ~n1527 & ~n11563;
  assign n11565 = ~n1550 & ~n1567;
  assign n11566 = ~n1563 & ~n11565;
  assign n11567 = ~n11564 & n11566;
  assign n11568 = n11564 & ~n11566;
  assign n11569 = ~n11567 & ~n11568;
  assign n11570 = ~n11562 & ~n11569;
  assign n11571 = ~n1753 & ~n11567;
  assign n11572 = ~n11568 & n11571;
  assign n11573 = ~n11561 & n11572;
  assign n11574 = ~n11570 & ~n11573;
  assign n11575 = n1758 & ~n1764;
  assign n11576 = ~n1768 & ~n11575;
  assign n11577 = ~n1439 & ~n1456;
  assign n11578 = ~n1452 & ~n11577;
  assign n11579 = ~n1475 & ~n1492;
  assign n11580 = ~n1488 & ~n11579;
  assign n11581 = ~n11578 & n11580;
  assign n11582 = n11578 & ~n11580;
  assign n11583 = ~n11581 & ~n11582;
  assign n11584 = ~n11576 & ~n11583;
  assign n11585 = ~n1768 & ~n11581;
  assign n11586 = ~n11582 & n11585;
  assign n11587 = ~n11575 & n11586;
  assign n11588 = ~n11584 & ~n11587;
  assign n11589 = ~n11574 & n11588;
  assign n11590 = n11574 & ~n11588;
  assign n11591 = ~n11589 & ~n11590;
  assign n11592 = ~n11560 & ~n11591;
  assign n11593 = n11560 & n11591;
  assign n11594 = ~n11592 & ~n11593;
  assign n11595 = ~n11558 & n11594;
  assign n11596 = n11558 & ~n11594;
  assign n11597 = ~n11595 & ~n11596;
  assign n11598 = ~n11522 & ~n11597;
  assign n11599 = n11522 & n11597;
  assign n11600 = ~n11598 & ~n11599;
  assign n11601 = ~n1202 & ~n1410;
  assign n11602 = ~n1412 & ~n11601;
  assign n11603 = ~n1195 & ~n1198;
  assign n11604 = ~n1199 & ~n11603;
  assign n11605 = n1178 & ~n1188;
  assign n11606 = ~n1192 & ~n11605;
  assign n11607 = ~n1112 & ~n1129;
  assign n11608 = ~n1125 & ~n11607;
  assign n11609 = ~n1148 & ~n1165;
  assign n11610 = ~n1161 & ~n11609;
  assign n11611 = ~n11608 & n11610;
  assign n11612 = n11608 & ~n11610;
  assign n11613 = ~n11611 & ~n11612;
  assign n11614 = ~n11606 & ~n11613;
  assign n11615 = ~n1192 & ~n11611;
  assign n11616 = ~n11612 & n11615;
  assign n11617 = ~n11605 & n11616;
  assign n11618 = ~n11614 & ~n11617;
  assign n11619 = n1038 & ~n1080;
  assign n11620 = ~n1084 & ~n11619;
  assign n11621 = ~n1070 & ~n1074;
  assign n11622 = ~n1066 & ~n11621;
  assign n11623 = ~n1030 & ~n1033;
  assign n11624 = ~n1036 & ~n11623;
  assign n11625 = ~n11622 & n11624;
  assign n11626 = n11622 & ~n11624;
  assign n11627 = ~n11625 & ~n11626;
  assign n11628 = ~n11620 & ~n11627;
  assign n11629 = ~n1084 & ~n11625;
  assign n11630 = ~n11626 & n11629;
  assign n11631 = ~n11619 & n11630;
  assign n11632 = ~n11628 & ~n11631;
  assign n11633 = ~n11618 & n11632;
  assign n11634 = n11618 & ~n11632;
  assign n11635 = ~n11633 & ~n11634;
  assign n11636 = ~n11604 & ~n11635;
  assign n11637 = n11604 & n11635;
  assign n11638 = ~n11636 & ~n11637;
  assign n11639 = ~n1291 & ~n1392;
  assign n11640 = ~n1394 & ~n11639;
  assign n11641 = n1238 & ~n1284;
  assign n11642 = ~n1288 & ~n11641;
  assign n11643 = ~n1270 & ~n1274;
  assign n11644 = ~n1266 & ~n11643;
  assign n11645 = ~n1230 & ~n1233;
  assign n11646 = ~n1236 & ~n11645;
  assign n11647 = ~n11644 & n11646;
  assign n11648 = n11644 & ~n11646;
  assign n11649 = ~n11647 & ~n11648;
  assign n11650 = ~n11642 & ~n11649;
  assign n11651 = ~n1288 & ~n11647;
  assign n11652 = ~n11648 & n11651;
  assign n11653 = ~n11641 & n11652;
  assign n11654 = ~n11650 & ~n11653;
  assign n11655 = n1327 & ~n1369;
  assign n11656 = ~n1373 & ~n11655;
  assign n11657 = ~n1359 & ~n1363;
  assign n11658 = ~n1355 & ~n11657;
  assign n11659 = ~n1319 & ~n1322;
  assign n11660 = ~n1325 & ~n11659;
  assign n11661 = ~n11658 & n11660;
  assign n11662 = n11658 & ~n11660;
  assign n11663 = ~n11661 & ~n11662;
  assign n11664 = ~n11656 & ~n11663;
  assign n11665 = ~n1373 & ~n11661;
  assign n11666 = ~n11662 & n11665;
  assign n11667 = ~n11655 & n11666;
  assign n11668 = ~n11664 & ~n11667;
  assign n11669 = ~n11654 & n11668;
  assign n11670 = n11654 & ~n11668;
  assign n11671 = ~n11669 & ~n11670;
  assign n11672 = ~n11640 & ~n11671;
  assign n11673 = n11640 & n11671;
  assign n11674 = ~n11672 & ~n11673;
  assign n11675 = ~n11638 & n11674;
  assign n11676 = n11638 & ~n11674;
  assign n11677 = ~n11675 & ~n11676;
  assign n11678 = ~n11602 & ~n11677;
  assign n11679 = n11602 & n11677;
  assign n11680 = ~n11678 & ~n11679;
  assign n11681 = ~n11600 & n11680;
  assign n11682 = n11600 & ~n11680;
  assign n11683 = ~n11681 & ~n11682;
  assign n11684 = ~n11520 & ~n11683;
  assign n11685 = n11520 & n11683;
  assign n11686 = ~n11684 & ~n11685;
  assign n11687 = ~n2274 & ~n2700;
  assign n11688 = ~n2702 & ~n11687;
  assign n11689 = ~n2267 & ~n2270;
  assign n11690 = ~n2271 & ~n11689;
  assign n11691 = ~n2260 & ~n2263;
  assign n11692 = ~n2264 & ~n11691;
  assign n11693 = n2243 & ~n2253;
  assign n11694 = ~n2257 & ~n11693;
  assign n11695 = ~n2150 & ~n2167;
  assign n11696 = ~n2163 & ~n11695;
  assign n11697 = ~n2186 & ~n2203;
  assign n11698 = ~n2199 & ~n11697;
  assign n11699 = ~n11696 & n11698;
  assign n11700 = n11696 & ~n11698;
  assign n11701 = ~n11699 & ~n11700;
  assign n11702 = ~n11694 & ~n11701;
  assign n11703 = ~n2257 & ~n11699;
  assign n11704 = ~n11700 & n11703;
  assign n11705 = ~n11693 & n11704;
  assign n11706 = ~n11702 & ~n11705;
  assign n11707 = n2219 & ~n2225;
  assign n11708 = ~n2229 & ~n11707;
  assign n11709 = ~n2075 & ~n2092;
  assign n11710 = ~n2088 & ~n11709;
  assign n11711 = ~n2111 & ~n2128;
  assign n11712 = ~n2124 & ~n11711;
  assign n11713 = ~n11710 & n11712;
  assign n11714 = n11710 & ~n11712;
  assign n11715 = ~n11713 & ~n11714;
  assign n11716 = ~n11708 & ~n11715;
  assign n11717 = ~n2229 & ~n11713;
  assign n11718 = ~n11714 & n11717;
  assign n11719 = ~n11707 & n11718;
  assign n11720 = ~n11716 & ~n11719;
  assign n11721 = ~n11706 & n11720;
  assign n11722 = n11706 & ~n11720;
  assign n11723 = ~n11721 & ~n11722;
  assign n11724 = ~n11692 & ~n11723;
  assign n11725 = n11692 & n11723;
  assign n11726 = ~n11724 & ~n11725;
  assign n11727 = ~n1945 & ~n2046;
  assign n11728 = ~n2048 & ~n11727;
  assign n11729 = n1892 & ~n1938;
  assign n11730 = ~n1942 & ~n11729;
  assign n11731 = ~n1924 & ~n1928;
  assign n11732 = ~n1920 & ~n11731;
  assign n11733 = ~n1884 & ~n1887;
  assign n11734 = ~n1890 & ~n11733;
  assign n11735 = ~n11732 & n11734;
  assign n11736 = n11732 & ~n11734;
  assign n11737 = ~n11735 & ~n11736;
  assign n11738 = ~n11730 & ~n11737;
  assign n11739 = ~n1942 & ~n11735;
  assign n11740 = ~n11736 & n11739;
  assign n11741 = ~n11729 & n11740;
  assign n11742 = ~n11738 & ~n11741;
  assign n11743 = n1981 & ~n2023;
  assign n11744 = ~n2027 & ~n11743;
  assign n11745 = ~n2013 & ~n2017;
  assign n11746 = ~n2009 & ~n11745;
  assign n11747 = ~n1973 & ~n1976;
  assign n11748 = ~n1979 & ~n11747;
  assign n11749 = ~n11746 & n11748;
  assign n11750 = n11746 & ~n11748;
  assign n11751 = ~n11749 & ~n11750;
  assign n11752 = ~n11744 & ~n11751;
  assign n11753 = ~n2027 & ~n11749;
  assign n11754 = ~n11750 & n11753;
  assign n11755 = ~n11743 & n11754;
  assign n11756 = ~n11752 & ~n11755;
  assign n11757 = ~n11742 & n11756;
  assign n11758 = n11742 & ~n11756;
  assign n11759 = ~n11757 & ~n11758;
  assign n11760 = ~n11728 & ~n11759;
  assign n11761 = n11728 & n11759;
  assign n11762 = ~n11760 & ~n11761;
  assign n11763 = ~n11726 & n11762;
  assign n11764 = n11726 & ~n11762;
  assign n11765 = ~n11763 & ~n11764;
  assign n11766 = ~n11690 & ~n11765;
  assign n11767 = n11690 & n11765;
  assign n11768 = ~n11766 & ~n11767;
  assign n11769 = ~n2474 & ~n2682;
  assign n11770 = ~n2684 & ~n11769;
  assign n11771 = ~n2467 & ~n2470;
  assign n11772 = ~n2471 & ~n11771;
  assign n11773 = n2450 & ~n2460;
  assign n11774 = ~n2464 & ~n11773;
  assign n11775 = ~n2384 & ~n2401;
  assign n11776 = ~n2397 & ~n11775;
  assign n11777 = ~n2420 & ~n2437;
  assign n11778 = ~n2433 & ~n11777;
  assign n11779 = ~n11776 & n11778;
  assign n11780 = n11776 & ~n11778;
  assign n11781 = ~n11779 & ~n11780;
  assign n11782 = ~n11774 & ~n11781;
  assign n11783 = ~n2464 & ~n11779;
  assign n11784 = ~n11780 & n11783;
  assign n11785 = ~n11773 & n11784;
  assign n11786 = ~n11782 & ~n11785;
  assign n11787 = n2310 & ~n2352;
  assign n11788 = ~n2356 & ~n11787;
  assign n11789 = ~n2342 & ~n2346;
  assign n11790 = ~n2338 & ~n11789;
  assign n11791 = ~n2302 & ~n2305;
  assign n11792 = ~n2308 & ~n11791;
  assign n11793 = ~n11790 & n11792;
  assign n11794 = n11790 & ~n11792;
  assign n11795 = ~n11793 & ~n11794;
  assign n11796 = ~n11788 & ~n11795;
  assign n11797 = ~n2356 & ~n11793;
  assign n11798 = ~n11794 & n11797;
  assign n11799 = ~n11787 & n11798;
  assign n11800 = ~n11796 & ~n11799;
  assign n11801 = ~n11786 & n11800;
  assign n11802 = n11786 & ~n11800;
  assign n11803 = ~n11801 & ~n11802;
  assign n11804 = ~n11772 & ~n11803;
  assign n11805 = n11772 & n11803;
  assign n11806 = ~n11804 & ~n11805;
  assign n11807 = ~n2563 & ~n2664;
  assign n11808 = ~n2666 & ~n11807;
  assign n11809 = n2510 & ~n2556;
  assign n11810 = ~n2560 & ~n11809;
  assign n11811 = ~n2542 & ~n2546;
  assign n11812 = ~n2538 & ~n11811;
  assign n11813 = ~n2502 & ~n2505;
  assign n11814 = ~n2508 & ~n11813;
  assign n11815 = ~n11812 & n11814;
  assign n11816 = n11812 & ~n11814;
  assign n11817 = ~n11815 & ~n11816;
  assign n11818 = ~n11810 & ~n11817;
  assign n11819 = ~n2560 & ~n11815;
  assign n11820 = ~n11816 & n11819;
  assign n11821 = ~n11809 & n11820;
  assign n11822 = ~n11818 & ~n11821;
  assign n11823 = n2599 & ~n2641;
  assign n11824 = ~n2645 & ~n11823;
  assign n11825 = ~n2631 & ~n2635;
  assign n11826 = ~n2627 & ~n11825;
  assign n11827 = ~n2591 & ~n2594;
  assign n11828 = ~n2597 & ~n11827;
  assign n11829 = ~n11826 & n11828;
  assign n11830 = n11826 & ~n11828;
  assign n11831 = ~n11829 & ~n11830;
  assign n11832 = ~n11824 & ~n11831;
  assign n11833 = ~n2645 & ~n11829;
  assign n11834 = ~n11830 & n11833;
  assign n11835 = ~n11823 & n11834;
  assign n11836 = ~n11832 & ~n11835;
  assign n11837 = ~n11822 & n11836;
  assign n11838 = n11822 & ~n11836;
  assign n11839 = ~n11837 & ~n11838;
  assign n11840 = ~n11808 & ~n11839;
  assign n11841 = n11808 & n11839;
  assign n11842 = ~n11840 & ~n11841;
  assign n11843 = ~n11806 & n11842;
  assign n11844 = n11806 & ~n11842;
  assign n11845 = ~n11843 & ~n11844;
  assign n11846 = ~n11770 & ~n11845;
  assign n11847 = n11770 & n11845;
  assign n11848 = ~n11846 & ~n11847;
  assign n11849 = ~n11768 & n11848;
  assign n11850 = n11768 & ~n11848;
  assign n11851 = ~n11849 & ~n11850;
  assign n11852 = ~n11688 & ~n11851;
  assign n11853 = n11688 & n11851;
  assign n11854 = ~n11852 & ~n11853;
  assign n11855 = ~n11686 & n11854;
  assign n11856 = n11686 & ~n11854;
  assign n11857 = ~n11855 & ~n11856;
  assign n11858 = ~n11518 & ~n11857;
  assign n11859 = n11518 & n11857;
  assign n11860 = ~n11858 & ~n11859;
  assign n11861 = ~n11516 & n11860;
  assign n11862 = n11516 & ~n11860;
  assign n11863 = ~n11861 & ~n11862;
  assign n11864 = ~n11172 & ~n11863;
  assign n11865 = n11172 & n11863;
  assign n11866 = ~n11864 & ~n11865;
  assign n11867 = ~n11170 & ~n11866;
  assign n11868 = ~n10047 & ~n11867;
  assign n11869 = ~n11168 & n11866;
  assign n11870 = ~n11169 & n11869;
  assign n11871 = ~n11868 & ~n11870;
  assign n11872 = ~n10468 & ~n11164;
  assign n11873 = ~n10049 & ~n11872;
  assign n11874 = n10468 & n11164;
  assign n11875 = ~n11873 & ~n11874;
  assign n11876 = ~n10814 & ~n11158;
  assign n11877 = ~n10470 & ~n11876;
  assign n11878 = n10814 & n11158;
  assign n11879 = ~n11877 & ~n11878;
  assign n11880 = ~n10984 & ~n11152;
  assign n11881 = ~n10816 & ~n11880;
  assign n11882 = n10984 & n11152;
  assign n11883 = ~n11881 & ~n11882;
  assign n11884 = ~n11066 & ~n11146;
  assign n11885 = ~n10986 & ~n11884;
  assign n11886 = n11066 & n11146;
  assign n11887 = ~n11885 & ~n11886;
  assign n11888 = ~n11104 & ~n11140;
  assign n11889 = ~n11068 & ~n11888;
  assign n11890 = n11104 & n11140;
  assign n11891 = ~n11889 & ~n11890;
  assign n11892 = ~n11120 & ~n11134;
  assign n11893 = ~n11106 & ~n11892;
  assign n11894 = ~n11119 & ~n11133;
  assign n11895 = ~n11130 & n11894;
  assign n11896 = ~n11116 & n11895;
  assign n11897 = ~n11893 & ~n11896;
  assign n11898 = ~n9915 & ~n11124;
  assign n11899 = ~n11121 & n11898;
  assign n11900 = n11126 & ~n11899;
  assign n11901 = ~n11122 & n11124;
  assign n11902 = ~n11900 & ~n11901;
  assign n11903 = ~n9830 & ~n11110;
  assign n11904 = ~n11107 & n11903;
  assign n11905 = n11112 & ~n11904;
  assign n11906 = ~n11108 & n11110;
  assign n11907 = ~n11905 & ~n11906;
  assign n11908 = ~n11902 & n11907;
  assign n11909 = n11902 & ~n11907;
  assign n11910 = ~n11908 & ~n11909;
  assign n11911 = ~n11897 & ~n11910;
  assign n11912 = ~n11896 & ~n11908;
  assign n11913 = ~n11909 & n11912;
  assign n11914 = ~n11893 & n11913;
  assign n11915 = ~n11911 & ~n11914;
  assign n11916 = ~n11084 & ~n11098;
  assign n11917 = ~n11070 & ~n11916;
  assign n11918 = ~n11083 & ~n11097;
  assign n11919 = ~n11094 & n11918;
  assign n11920 = ~n11080 & n11919;
  assign n11921 = ~n11917 & ~n11920;
  assign n11922 = ~n9626 & ~n11088;
  assign n11923 = ~n11085 & n11922;
  assign n11924 = n11090 & ~n11923;
  assign n11925 = ~n11086 & n11088;
  assign n11926 = ~n11924 & ~n11925;
  assign n11927 = ~n9734 & ~n11074;
  assign n11928 = ~n11071 & n11927;
  assign n11929 = n11076 & ~n11928;
  assign n11930 = ~n11072 & n11074;
  assign n11931 = ~n11929 & ~n11930;
  assign n11932 = ~n11926 & n11931;
  assign n11933 = n11926 & ~n11931;
  assign n11934 = ~n11932 & ~n11933;
  assign n11935 = ~n11921 & ~n11934;
  assign n11936 = ~n11920 & ~n11932;
  assign n11937 = ~n11933 & n11936;
  assign n11938 = ~n11917 & n11937;
  assign n11939 = ~n11935 & ~n11938;
  assign n11940 = ~n11915 & n11939;
  assign n11941 = n11915 & ~n11939;
  assign n11942 = ~n11940 & ~n11941;
  assign n11943 = ~n11891 & ~n11942;
  assign n11944 = n11891 & n11942;
  assign n11945 = ~n11943 & ~n11944;
  assign n11946 = ~n11024 & ~n11060;
  assign n11947 = ~n10988 & ~n11946;
  assign n11948 = n11024 & n11060;
  assign n11949 = ~n11947 & ~n11948;
  assign n11950 = ~n11040 & ~n11054;
  assign n11951 = ~n11026 & ~n11950;
  assign n11952 = ~n11039 & ~n11053;
  assign n11953 = ~n11050 & n11952;
  assign n11954 = ~n11036 & n11953;
  assign n11955 = ~n11951 & ~n11954;
  assign n11956 = ~n9297 & ~n11044;
  assign n11957 = ~n11041 & n11956;
  assign n11958 = n11046 & ~n11957;
  assign n11959 = ~n11042 & n11044;
  assign n11960 = ~n11958 & ~n11959;
  assign n11961 = ~n9212 & ~n11030;
  assign n11962 = ~n11027 & n11961;
  assign n11963 = n11032 & ~n11962;
  assign n11964 = ~n11028 & n11030;
  assign n11965 = ~n11963 & ~n11964;
  assign n11966 = ~n11960 & n11965;
  assign n11967 = n11960 & ~n11965;
  assign n11968 = ~n11966 & ~n11967;
  assign n11969 = ~n11955 & ~n11968;
  assign n11970 = ~n11954 & ~n11966;
  assign n11971 = ~n11967 & n11970;
  assign n11972 = ~n11951 & n11971;
  assign n11973 = ~n11969 & ~n11972;
  assign n11974 = ~n11004 & ~n11018;
  assign n11975 = ~n10990 & ~n11974;
  assign n11976 = ~n11003 & ~n11017;
  assign n11977 = ~n11014 & n11976;
  assign n11978 = ~n11000 & n11977;
  assign n11979 = ~n11975 & ~n11978;
  assign n11980 = ~n9499 & ~n11008;
  assign n11981 = ~n11005 & n11980;
  assign n11982 = n11010 & ~n11981;
  assign n11983 = ~n11006 & n11008;
  assign n11984 = ~n11982 & ~n11983;
  assign n11985 = ~n9527 & ~n10994;
  assign n11986 = ~n10991 & n11985;
  assign n11987 = n10996 & ~n11986;
  assign n11988 = ~n10992 & n10994;
  assign n11989 = ~n11987 & ~n11988;
  assign n11990 = ~n11984 & n11989;
  assign n11991 = n11984 & ~n11989;
  assign n11992 = ~n11990 & ~n11991;
  assign n11993 = ~n11979 & ~n11992;
  assign n11994 = ~n11978 & ~n11990;
  assign n11995 = ~n11991 & n11994;
  assign n11996 = ~n11975 & n11995;
  assign n11997 = ~n11993 & ~n11996;
  assign n11998 = ~n11973 & n11997;
  assign n11999 = n11973 & ~n11997;
  assign n12000 = ~n11998 & ~n11999;
  assign n12001 = ~n11949 & ~n12000;
  assign n12002 = n11949 & n12000;
  assign n12003 = ~n12001 & ~n12002;
  assign n12004 = ~n11945 & n12003;
  assign n12005 = n11945 & ~n12003;
  assign n12006 = ~n12004 & ~n12005;
  assign n12007 = ~n11887 & ~n12006;
  assign n12008 = n11887 & n12006;
  assign n12009 = ~n12007 & ~n12008;
  assign n12010 = ~n10898 & ~n10978;
  assign n12011 = ~n10818 & ~n12010;
  assign n12012 = n10898 & n10978;
  assign n12013 = ~n12011 & ~n12012;
  assign n12014 = ~n10936 & ~n10972;
  assign n12015 = ~n10900 & ~n12014;
  assign n12016 = n10936 & n10972;
  assign n12017 = ~n12015 & ~n12016;
  assign n12018 = ~n10952 & ~n10966;
  assign n12019 = ~n10938 & ~n12018;
  assign n12020 = ~n10951 & ~n10965;
  assign n12021 = ~n10962 & n12020;
  assign n12022 = ~n10948 & n12021;
  assign n12023 = ~n12019 & ~n12022;
  assign n12024 = ~n8643 & ~n10956;
  assign n12025 = ~n10953 & n12024;
  assign n12026 = n10958 & ~n12025;
  assign n12027 = ~n10954 & n10956;
  assign n12028 = ~n12026 & ~n12027;
  assign n12029 = ~n8558 & ~n10942;
  assign n12030 = ~n10939 & n12029;
  assign n12031 = n10944 & ~n12030;
  assign n12032 = ~n10940 & n10942;
  assign n12033 = ~n12031 & ~n12032;
  assign n12034 = ~n12028 & n12033;
  assign n12035 = n12028 & ~n12033;
  assign n12036 = ~n12034 & ~n12035;
  assign n12037 = ~n12023 & ~n12036;
  assign n12038 = ~n12022 & ~n12034;
  assign n12039 = ~n12035 & n12038;
  assign n12040 = ~n12019 & n12039;
  assign n12041 = ~n12037 & ~n12040;
  assign n12042 = ~n10916 & ~n10930;
  assign n12043 = ~n10902 & ~n12042;
  assign n12044 = ~n10915 & ~n10929;
  assign n12045 = ~n10926 & n12044;
  assign n12046 = ~n10912 & n12045;
  assign n12047 = ~n12043 & ~n12046;
  assign n12048 = ~n8354 & ~n10920;
  assign n12049 = ~n10917 & n12048;
  assign n12050 = n10922 & ~n12049;
  assign n12051 = ~n10918 & n10920;
  assign n12052 = ~n12050 & ~n12051;
  assign n12053 = ~n8462 & ~n10906;
  assign n12054 = ~n10903 & n12053;
  assign n12055 = n10908 & ~n12054;
  assign n12056 = ~n10904 & n10906;
  assign n12057 = ~n12055 & ~n12056;
  assign n12058 = ~n12052 & n12057;
  assign n12059 = n12052 & ~n12057;
  assign n12060 = ~n12058 & ~n12059;
  assign n12061 = ~n12047 & ~n12060;
  assign n12062 = ~n12046 & ~n12058;
  assign n12063 = ~n12059 & n12062;
  assign n12064 = ~n12043 & n12063;
  assign n12065 = ~n12061 & ~n12064;
  assign n12066 = ~n12041 & n12065;
  assign n12067 = n12041 & ~n12065;
  assign n12068 = ~n12066 & ~n12067;
  assign n12069 = ~n12017 & ~n12068;
  assign n12070 = n12017 & n12068;
  assign n12071 = ~n12069 & ~n12070;
  assign n12072 = ~n10856 & ~n10892;
  assign n12073 = ~n10820 & ~n12072;
  assign n12074 = n10856 & n10892;
  assign n12075 = ~n12073 & ~n12074;
  assign n12076 = ~n10872 & ~n10886;
  assign n12077 = ~n10858 & ~n12076;
  assign n12078 = ~n10871 & ~n10885;
  assign n12079 = ~n10882 & n12078;
  assign n12080 = ~n10868 & n12079;
  assign n12081 = ~n12077 & ~n12080;
  assign n12082 = ~n9038 & ~n10876;
  assign n12083 = ~n10873 & n12082;
  assign n12084 = n10878 & ~n12083;
  assign n12085 = ~n10874 & n10876;
  assign n12086 = ~n12084 & ~n12085;
  assign n12087 = ~n9023 & ~n10862;
  assign n12088 = ~n10859 & n12087;
  assign n12089 = n10864 & ~n12088;
  assign n12090 = ~n10860 & n10862;
  assign n12091 = ~n12089 & ~n12090;
  assign n12092 = ~n12086 & n12091;
  assign n12093 = n12086 & ~n12091;
  assign n12094 = ~n12092 & ~n12093;
  assign n12095 = ~n12081 & ~n12094;
  assign n12096 = ~n12080 & ~n12092;
  assign n12097 = ~n12093 & n12096;
  assign n12098 = ~n12077 & n12097;
  assign n12099 = ~n12095 & ~n12098;
  assign n12100 = ~n10836 & ~n10850;
  assign n12101 = ~n10822 & ~n12100;
  assign n12102 = ~n10835 & ~n10849;
  assign n12103 = ~n10846 & n12102;
  assign n12104 = ~n10832 & n12103;
  assign n12105 = ~n12101 & ~n12104;
  assign n12106 = ~n9074 & ~n10840;
  assign n12107 = ~n10837 & n12106;
  assign n12108 = n10842 & ~n12107;
  assign n12109 = ~n10838 & n10840;
  assign n12110 = ~n12108 & ~n12109;
  assign n12111 = ~n9102 & ~n10826;
  assign n12112 = ~n10823 & n12111;
  assign n12113 = n10828 & ~n12112;
  assign n12114 = ~n10824 & n10826;
  assign n12115 = ~n12113 & ~n12114;
  assign n12116 = ~n12110 & n12115;
  assign n12117 = n12110 & ~n12115;
  assign n12118 = ~n12116 & ~n12117;
  assign n12119 = ~n12105 & ~n12118;
  assign n12120 = ~n12104 & ~n12116;
  assign n12121 = ~n12117 & n12120;
  assign n12122 = ~n12101 & n12121;
  assign n12123 = ~n12119 & ~n12122;
  assign n12124 = ~n12099 & n12123;
  assign n12125 = n12099 & ~n12123;
  assign n12126 = ~n12124 & ~n12125;
  assign n12127 = ~n12075 & ~n12126;
  assign n12128 = n12075 & n12126;
  assign n12129 = ~n12127 & ~n12128;
  assign n12130 = ~n12071 & n12129;
  assign n12131 = n12071 & ~n12129;
  assign n12132 = ~n12130 & ~n12131;
  assign n12133 = ~n12013 & ~n12132;
  assign n12134 = n12013 & n12132;
  assign n12135 = ~n12133 & ~n12134;
  assign n12136 = ~n12009 & n12135;
  assign n12137 = n12009 & ~n12135;
  assign n12138 = ~n12136 & ~n12137;
  assign n12139 = ~n11883 & ~n12138;
  assign n12140 = n11883 & n12138;
  assign n12141 = ~n12139 & ~n12140;
  assign n12142 = ~n10640 & ~n10808;
  assign n12143 = ~n10472 & ~n12142;
  assign n12144 = n10640 & n10808;
  assign n12145 = ~n12143 & ~n12144;
  assign n12146 = ~n10722 & ~n10802;
  assign n12147 = ~n10642 & ~n12146;
  assign n12148 = n10722 & n10802;
  assign n12149 = ~n12147 & ~n12148;
  assign n12150 = ~n10760 & ~n10796;
  assign n12151 = ~n10724 & ~n12150;
  assign n12152 = n10760 & n10796;
  assign n12153 = ~n12151 & ~n12152;
  assign n12154 = ~n10776 & ~n10790;
  assign n12155 = ~n10762 & ~n12154;
  assign n12156 = ~n10775 & ~n10789;
  assign n12157 = ~n10786 & n12156;
  assign n12158 = ~n10772 & n12157;
  assign n12159 = ~n12155 & ~n12158;
  assign n12160 = ~n7335 & ~n10780;
  assign n12161 = ~n10777 & n12160;
  assign n12162 = n10782 & ~n12161;
  assign n12163 = ~n10778 & n10780;
  assign n12164 = ~n12162 & ~n12163;
  assign n12165 = ~n7250 & ~n10766;
  assign n12166 = ~n10763 & n12165;
  assign n12167 = n10768 & ~n12166;
  assign n12168 = ~n10764 & n10766;
  assign n12169 = ~n12167 & ~n12168;
  assign n12170 = ~n12164 & n12169;
  assign n12171 = n12164 & ~n12169;
  assign n12172 = ~n12170 & ~n12171;
  assign n12173 = ~n12159 & ~n12172;
  assign n12174 = ~n12158 & ~n12170;
  assign n12175 = ~n12171 & n12174;
  assign n12176 = ~n12155 & n12175;
  assign n12177 = ~n12173 & ~n12176;
  assign n12178 = ~n10740 & ~n10754;
  assign n12179 = ~n10726 & ~n12178;
  assign n12180 = ~n10739 & ~n10753;
  assign n12181 = ~n10750 & n12180;
  assign n12182 = ~n10736 & n12181;
  assign n12183 = ~n12179 & ~n12182;
  assign n12184 = ~n7046 & ~n10744;
  assign n12185 = ~n10741 & n12184;
  assign n12186 = n10746 & ~n12185;
  assign n12187 = ~n10742 & n10744;
  assign n12188 = ~n12186 & ~n12187;
  assign n12189 = ~n7154 & ~n10730;
  assign n12190 = ~n10727 & n12189;
  assign n12191 = n10732 & ~n12190;
  assign n12192 = ~n10728 & n10730;
  assign n12193 = ~n12191 & ~n12192;
  assign n12194 = ~n12188 & n12193;
  assign n12195 = n12188 & ~n12193;
  assign n12196 = ~n12194 & ~n12195;
  assign n12197 = ~n12183 & ~n12196;
  assign n12198 = ~n12182 & ~n12194;
  assign n12199 = ~n12195 & n12198;
  assign n12200 = ~n12179 & n12199;
  assign n12201 = ~n12197 & ~n12200;
  assign n12202 = ~n12177 & n12201;
  assign n12203 = n12177 & ~n12201;
  assign n12204 = ~n12202 & ~n12203;
  assign n12205 = ~n12153 & ~n12204;
  assign n12206 = n12153 & n12204;
  assign n12207 = ~n12205 & ~n12206;
  assign n12208 = ~n10680 & ~n10716;
  assign n12209 = ~n10644 & ~n12208;
  assign n12210 = n10680 & n10716;
  assign n12211 = ~n12209 & ~n12210;
  assign n12212 = ~n10696 & ~n10710;
  assign n12213 = ~n10682 & ~n12212;
  assign n12214 = ~n10695 & ~n10709;
  assign n12215 = ~n10706 & n12214;
  assign n12216 = ~n10692 & n12215;
  assign n12217 = ~n12213 & ~n12216;
  assign n12218 = ~n6717 & ~n10700;
  assign n12219 = ~n10697 & n12218;
  assign n12220 = n10702 & ~n12219;
  assign n12221 = ~n10698 & n10700;
  assign n12222 = ~n12220 & ~n12221;
  assign n12223 = ~n6632 & ~n10686;
  assign n12224 = ~n10683 & n12223;
  assign n12225 = n10688 & ~n12224;
  assign n12226 = ~n10684 & n10686;
  assign n12227 = ~n12225 & ~n12226;
  assign n12228 = ~n12222 & n12227;
  assign n12229 = n12222 & ~n12227;
  assign n12230 = ~n12228 & ~n12229;
  assign n12231 = ~n12217 & ~n12230;
  assign n12232 = ~n12216 & ~n12228;
  assign n12233 = ~n12229 & n12232;
  assign n12234 = ~n12213 & n12233;
  assign n12235 = ~n12231 & ~n12234;
  assign n12236 = ~n10660 & ~n10674;
  assign n12237 = ~n10646 & ~n12236;
  assign n12238 = ~n10659 & ~n10673;
  assign n12239 = ~n10670 & n12238;
  assign n12240 = ~n10656 & n12239;
  assign n12241 = ~n12237 & ~n12240;
  assign n12242 = ~n6919 & ~n10664;
  assign n12243 = ~n10661 & n12242;
  assign n12244 = n10666 & ~n12243;
  assign n12245 = ~n10662 & n10664;
  assign n12246 = ~n12244 & ~n12245;
  assign n12247 = ~n6947 & ~n10650;
  assign n12248 = ~n10647 & n12247;
  assign n12249 = n10652 & ~n12248;
  assign n12250 = ~n10648 & n10650;
  assign n12251 = ~n12249 & ~n12250;
  assign n12252 = ~n12246 & n12251;
  assign n12253 = n12246 & ~n12251;
  assign n12254 = ~n12252 & ~n12253;
  assign n12255 = ~n12241 & ~n12254;
  assign n12256 = ~n12240 & ~n12252;
  assign n12257 = ~n12253 & n12256;
  assign n12258 = ~n12237 & n12257;
  assign n12259 = ~n12255 & ~n12258;
  assign n12260 = ~n12235 & n12259;
  assign n12261 = n12235 & ~n12259;
  assign n12262 = ~n12260 & ~n12261;
  assign n12263 = ~n12211 & ~n12262;
  assign n12264 = n12211 & n12262;
  assign n12265 = ~n12263 & ~n12264;
  assign n12266 = ~n12207 & n12265;
  assign n12267 = n12207 & ~n12265;
  assign n12268 = ~n12266 & ~n12267;
  assign n12269 = ~n12149 & ~n12268;
  assign n12270 = n12149 & n12268;
  assign n12271 = ~n12269 & ~n12270;
  assign n12272 = ~n10554 & ~n10634;
  assign n12273 = ~n10474 & ~n12272;
  assign n12274 = n10554 & n10634;
  assign n12275 = ~n12273 & ~n12274;
  assign n12276 = ~n10592 & ~n10628;
  assign n12277 = ~n10556 & ~n12276;
  assign n12278 = n10592 & n10628;
  assign n12279 = ~n12277 & ~n12278;
  assign n12280 = ~n10608 & ~n10622;
  assign n12281 = ~n10594 & ~n12280;
  assign n12282 = ~n10607 & ~n10621;
  assign n12283 = ~n10618 & n12282;
  assign n12284 = ~n10604 & n12283;
  assign n12285 = ~n12281 & ~n12284;
  assign n12286 = ~n8110 & ~n10612;
  assign n12287 = ~n10609 & n12286;
  assign n12288 = n10614 & ~n12287;
  assign n12289 = ~n10610 & n10612;
  assign n12290 = ~n12288 & ~n12289;
  assign n12291 = ~n8095 & ~n10598;
  assign n12292 = ~n10595 & n12291;
  assign n12293 = n10600 & ~n12292;
  assign n12294 = ~n10596 & n10598;
  assign n12295 = ~n12293 & ~n12294;
  assign n12296 = ~n12290 & n12295;
  assign n12297 = n12290 & ~n12295;
  assign n12298 = ~n12296 & ~n12297;
  assign n12299 = ~n12285 & ~n12298;
  assign n12300 = ~n12284 & ~n12296;
  assign n12301 = ~n12297 & n12300;
  assign n12302 = ~n12281 & n12301;
  assign n12303 = ~n12299 & ~n12302;
  assign n12304 = ~n10572 & ~n10586;
  assign n12305 = ~n10558 & ~n12304;
  assign n12306 = ~n10571 & ~n10585;
  assign n12307 = ~n10582 & n12306;
  assign n12308 = ~n10568 & n12307;
  assign n12309 = ~n12305 & ~n12308;
  assign n12310 = ~n8041 & ~n10576;
  assign n12311 = ~n10573 & n12310;
  assign n12312 = n10578 & ~n12311;
  assign n12313 = ~n10574 & n10576;
  assign n12314 = ~n12312 & ~n12313;
  assign n12315 = ~n8069 & ~n10562;
  assign n12316 = ~n10559 & n12315;
  assign n12317 = n10564 & ~n12316;
  assign n12318 = ~n10560 & n10562;
  assign n12319 = ~n12317 & ~n12318;
  assign n12320 = ~n12314 & n12319;
  assign n12321 = n12314 & ~n12319;
  assign n12322 = ~n12320 & ~n12321;
  assign n12323 = ~n12309 & ~n12322;
  assign n12324 = ~n12308 & ~n12320;
  assign n12325 = ~n12321 & n12324;
  assign n12326 = ~n12305 & n12325;
  assign n12327 = ~n12323 & ~n12326;
  assign n12328 = ~n12303 & n12327;
  assign n12329 = n12303 & ~n12327;
  assign n12330 = ~n12328 & ~n12329;
  assign n12331 = ~n12279 & ~n12330;
  assign n12332 = n12279 & n12330;
  assign n12333 = ~n12331 & ~n12332;
  assign n12334 = ~n10512 & ~n10548;
  assign n12335 = ~n10476 & ~n12334;
  assign n12336 = n10512 & n10548;
  assign n12337 = ~n12335 & ~n12336;
  assign n12338 = ~n10528 & ~n10542;
  assign n12339 = ~n10514 & ~n12338;
  assign n12340 = ~n10527 & ~n10541;
  assign n12341 = ~n10538 & n12340;
  assign n12342 = ~n10524 & n12341;
  assign n12343 = ~n12339 & ~n12342;
  assign n12344 = ~n8177 & ~n10532;
  assign n12345 = ~n10529 & n12344;
  assign n12346 = n10534 & ~n12345;
  assign n12347 = ~n10530 & n10532;
  assign n12348 = ~n12346 & ~n12347;
  assign n12349 = ~n8162 & ~n10518;
  assign n12350 = ~n10515 & n12349;
  assign n12351 = n10520 & ~n12350;
  assign n12352 = ~n10516 & n10518;
  assign n12353 = ~n12351 & ~n12352;
  assign n12354 = ~n12348 & n12353;
  assign n12355 = n12348 & ~n12353;
  assign n12356 = ~n12354 & ~n12355;
  assign n12357 = ~n12343 & ~n12356;
  assign n12358 = ~n12342 & ~n12354;
  assign n12359 = ~n12355 & n12358;
  assign n12360 = ~n12339 & n12359;
  assign n12361 = ~n12357 & ~n12360;
  assign n12362 = ~n10492 & ~n10506;
  assign n12363 = ~n10478 & ~n12362;
  assign n12364 = ~n10491 & ~n10505;
  assign n12365 = ~n10502 & n12364;
  assign n12366 = ~n10488 & n12365;
  assign n12367 = ~n12363 & ~n12366;
  assign n12368 = ~n8213 & ~n10496;
  assign n12369 = ~n10493 & n12368;
  assign n12370 = n10498 & ~n12369;
  assign n12371 = ~n10494 & n10496;
  assign n12372 = ~n12370 & ~n12371;
  assign n12373 = ~n8241 & ~n10482;
  assign n12374 = ~n10479 & n12373;
  assign n12375 = n10484 & ~n12374;
  assign n12376 = ~n10480 & n10482;
  assign n12377 = ~n12375 & ~n12376;
  assign n12378 = ~n12372 & n12377;
  assign n12379 = n12372 & ~n12377;
  assign n12380 = ~n12378 & ~n12379;
  assign n12381 = ~n12367 & ~n12380;
  assign n12382 = ~n12366 & ~n12378;
  assign n12383 = ~n12379 & n12382;
  assign n12384 = ~n12363 & n12383;
  assign n12385 = ~n12381 & ~n12384;
  assign n12386 = ~n12361 & n12385;
  assign n12387 = n12361 & ~n12385;
  assign n12388 = ~n12386 & ~n12387;
  assign n12389 = ~n12337 & ~n12388;
  assign n12390 = n12337 & n12388;
  assign n12391 = ~n12389 & ~n12390;
  assign n12392 = ~n12333 & n12391;
  assign n12393 = n12333 & ~n12391;
  assign n12394 = ~n12392 & ~n12393;
  assign n12395 = ~n12275 & ~n12394;
  assign n12396 = n12275 & n12394;
  assign n12397 = ~n12395 & ~n12396;
  assign n12398 = ~n12271 & n12397;
  assign n12399 = n12271 & ~n12397;
  assign n12400 = ~n12398 & ~n12399;
  assign n12401 = ~n12145 & ~n12400;
  assign n12402 = n12145 & n12400;
  assign n12403 = ~n12401 & ~n12402;
  assign n12404 = ~n12141 & n12403;
  assign n12405 = n12141 & ~n12403;
  assign n12406 = ~n12404 & ~n12405;
  assign n12407 = ~n11879 & ~n12406;
  assign n12408 = n11879 & n12406;
  assign n12409 = ~n12407 & ~n12408;
  assign n12410 = ~n10460 & ~n10463;
  assign n12411 = ~n10051 & ~n12410;
  assign n12412 = ~n10292 & n10460;
  assign n12413 = ~n10291 & n12412;
  assign n12414 = ~n12411 & ~n12413;
  assign n12415 = ~n10285 & ~n10288;
  assign n12416 = ~n10053 & ~n12415;
  assign n12417 = ~n10205 & n10285;
  assign n12418 = ~n10204 & n12417;
  assign n12419 = ~n12416 & ~n12418;
  assign n12420 = ~n10120 & ~n10200;
  assign n12421 = ~n10055 & ~n12420;
  assign n12422 = n10120 & n10200;
  assign n12423 = ~n12421 & ~n12422;
  assign n12424 = ~n10158 & ~n10194;
  assign n12425 = ~n10122 & ~n12424;
  assign n12426 = n10158 & n10194;
  assign n12427 = ~n12425 & ~n12426;
  assign n12428 = ~n10174 & ~n10188;
  assign n12429 = ~n10160 & ~n12428;
  assign n12430 = ~n10173 & ~n10187;
  assign n12431 = ~n10184 & n12430;
  assign n12432 = ~n10170 & n12431;
  assign n12433 = ~n12429 & ~n12432;
  assign n12434 = ~n5589 & ~n10178;
  assign n12435 = ~n10175 & n12434;
  assign n12436 = n10180 & ~n12435;
  assign n12437 = ~n10176 & n10178;
  assign n12438 = ~n12436 & ~n12437;
  assign n12439 = ~n5504 & ~n10164;
  assign n12440 = ~n10161 & n12439;
  assign n12441 = n10166 & ~n12440;
  assign n12442 = ~n10162 & n10164;
  assign n12443 = ~n12441 & ~n12442;
  assign n12444 = ~n12438 & n12443;
  assign n12445 = n12438 & ~n12443;
  assign n12446 = ~n12444 & ~n12445;
  assign n12447 = ~n12433 & ~n12446;
  assign n12448 = ~n12432 & ~n12444;
  assign n12449 = ~n12445 & n12448;
  assign n12450 = ~n12429 & n12449;
  assign n12451 = ~n12447 & ~n12450;
  assign n12452 = ~n10138 & ~n10152;
  assign n12453 = ~n10124 & ~n12452;
  assign n12454 = ~n10137 & ~n10151;
  assign n12455 = ~n10148 & n12454;
  assign n12456 = ~n10134 & n12455;
  assign n12457 = ~n12453 & ~n12456;
  assign n12458 = ~n5300 & ~n10142;
  assign n12459 = ~n10139 & n12458;
  assign n12460 = n10144 & ~n12459;
  assign n12461 = ~n10140 & n10142;
  assign n12462 = ~n12460 & ~n12461;
  assign n12463 = ~n5408 & ~n10128;
  assign n12464 = ~n10125 & n12463;
  assign n12465 = n10130 & ~n12464;
  assign n12466 = ~n10126 & n10128;
  assign n12467 = ~n12465 & ~n12466;
  assign n12468 = ~n12462 & n12467;
  assign n12469 = n12462 & ~n12467;
  assign n12470 = ~n12468 & ~n12469;
  assign n12471 = ~n12457 & ~n12470;
  assign n12472 = ~n12456 & ~n12468;
  assign n12473 = ~n12469 & n12472;
  assign n12474 = ~n12453 & n12473;
  assign n12475 = ~n12471 & ~n12474;
  assign n12476 = ~n12451 & n12475;
  assign n12477 = n12451 & ~n12475;
  assign n12478 = ~n12476 & ~n12477;
  assign n12479 = ~n12427 & ~n12478;
  assign n12480 = n12427 & n12478;
  assign n12481 = ~n12479 & ~n12480;
  assign n12482 = ~n10078 & ~n10114;
  assign n12483 = ~n10057 & ~n12482;
  assign n12484 = n10078 & ~n10112;
  assign n12485 = ~n10113 & n12484;
  assign n12486 = ~n12483 & ~n12485;
  assign n12487 = ~n5208 & n10071;
  assign n12488 = ~n10058 & n12487;
  assign n12489 = n10068 & ~n12488;
  assign n12490 = ~n10059 & ~n10071;
  assign n12491 = ~n12489 & ~n12490;
  assign n12492 = ~n10061 & ~n10063;
  assign n12493 = ~n12491 & n12492;
  assign n12494 = ~n12489 & ~n12492;
  assign n12495 = ~n12490 & n12494;
  assign n12496 = ~n12493 & ~n12495;
  assign n12497 = ~n10094 & ~n10108;
  assign n12498 = ~n10080 & ~n12497;
  assign n12499 = ~n10093 & ~n10107;
  assign n12500 = ~n10104 & n12499;
  assign n12501 = ~n10090 & n12500;
  assign n12502 = ~n12498 & ~n12501;
  assign n12503 = ~n5061 & ~n10098;
  assign n12504 = ~n10095 & n12503;
  assign n12505 = n10100 & ~n12504;
  assign n12506 = ~n10096 & n10098;
  assign n12507 = ~n12505 & ~n12506;
  assign n12508 = ~n4976 & ~n10084;
  assign n12509 = ~n10081 & n12508;
  assign n12510 = n10086 & ~n12509;
  assign n12511 = ~n10082 & n10084;
  assign n12512 = ~n12510 & ~n12511;
  assign n12513 = ~n12507 & n12512;
  assign n12514 = n12507 & ~n12512;
  assign n12515 = ~n12513 & ~n12514;
  assign n12516 = ~n12502 & ~n12515;
  assign n12517 = ~n12501 & ~n12513;
  assign n12518 = ~n12514 & n12517;
  assign n12519 = ~n12498 & n12518;
  assign n12520 = ~n12516 & ~n12519;
  assign n12521 = ~n12496 & ~n12520;
  assign n12522 = n12496 & n12520;
  assign n12523 = ~n12521 & ~n12522;
  assign n12524 = ~n12486 & n12523;
  assign n12525 = n12486 & ~n12523;
  assign n12526 = ~n12524 & ~n12525;
  assign n12527 = ~n12481 & n12526;
  assign n12528 = n12481 & ~n12526;
  assign n12529 = ~n12527 & ~n12528;
  assign n12530 = ~n12423 & ~n12529;
  assign n12531 = n12423 & n12529;
  assign n12532 = ~n12530 & ~n12531;
  assign n12533 = ~n10243 & ~n10279;
  assign n12534 = ~n10207 & ~n12533;
  assign n12535 = n10243 & n10279;
  assign n12536 = ~n12534 & ~n12535;
  assign n12537 = ~n10259 & ~n10273;
  assign n12538 = ~n10245 & ~n12537;
  assign n12539 = ~n10258 & ~n10272;
  assign n12540 = ~n10269 & n12539;
  assign n12541 = ~n10255 & n12540;
  assign n12542 = ~n12538 & ~n12541;
  assign n12543 = ~n4643 & ~n10263;
  assign n12544 = ~n10260 & n12543;
  assign n12545 = n10265 & ~n12544;
  assign n12546 = ~n10261 & n10263;
  assign n12547 = ~n12545 & ~n12546;
  assign n12548 = ~n4558 & ~n10249;
  assign n12549 = ~n10246 & n12548;
  assign n12550 = n10251 & ~n12549;
  assign n12551 = ~n10247 & n10249;
  assign n12552 = ~n12550 & ~n12551;
  assign n12553 = ~n12547 & n12552;
  assign n12554 = n12547 & ~n12552;
  assign n12555 = ~n12553 & ~n12554;
  assign n12556 = ~n12542 & ~n12555;
  assign n12557 = ~n12541 & ~n12553;
  assign n12558 = ~n12554 & n12557;
  assign n12559 = ~n12538 & n12558;
  assign n12560 = ~n12556 & ~n12559;
  assign n12561 = ~n10223 & ~n10237;
  assign n12562 = ~n10209 & ~n12561;
  assign n12563 = ~n10222 & ~n10236;
  assign n12564 = ~n10233 & n12563;
  assign n12565 = ~n10219 & n12564;
  assign n12566 = ~n12562 & ~n12565;
  assign n12567 = ~n4845 & ~n10227;
  assign n12568 = ~n10224 & n12567;
  assign n12569 = n10229 & ~n12568;
  assign n12570 = ~n10225 & n10227;
  assign n12571 = ~n12569 & ~n12570;
  assign n12572 = ~n4873 & ~n10213;
  assign n12573 = ~n10210 & n12572;
  assign n12574 = n10215 & ~n12573;
  assign n12575 = ~n10211 & n10213;
  assign n12576 = ~n12574 & ~n12575;
  assign n12577 = ~n12571 & n12576;
  assign n12578 = n12571 & ~n12576;
  assign n12579 = ~n12577 & ~n12578;
  assign n12580 = ~n12566 & ~n12579;
  assign n12581 = ~n12565 & ~n12577;
  assign n12582 = ~n12578 & n12581;
  assign n12583 = ~n12562 & n12582;
  assign n12584 = ~n12580 & ~n12583;
  assign n12585 = ~n12560 & n12584;
  assign n12586 = n12560 & ~n12584;
  assign n12587 = ~n12585 & ~n12586;
  assign n12588 = ~n12536 & ~n12587;
  assign n12589 = n12536 & n12587;
  assign n12590 = ~n12588 & ~n12589;
  assign n12591 = ~n12532 & n12590;
  assign n12592 = ~n12530 & ~n12590;
  assign n12593 = ~n12531 & n12592;
  assign n12594 = ~n12591 & ~n12593;
  assign n12595 = ~n12419 & ~n12594;
  assign n12596 = n12419 & n12594;
  assign n12597 = ~n12595 & ~n12596;
  assign n12598 = ~n10374 & ~n10454;
  assign n12599 = ~n10294 & ~n12598;
  assign n12600 = n10374 & n10454;
  assign n12601 = ~n12599 & ~n12600;
  assign n12602 = ~n10412 & ~n10448;
  assign n12603 = ~n10376 & ~n12602;
  assign n12604 = n10412 & n10448;
  assign n12605 = ~n12603 & ~n12604;
  assign n12606 = ~n10428 & ~n10442;
  assign n12607 = ~n10414 & ~n12606;
  assign n12608 = ~n10427 & ~n10441;
  assign n12609 = ~n10438 & n12608;
  assign n12610 = ~n10424 & n12609;
  assign n12611 = ~n12607 & ~n12610;
  assign n12612 = ~n6384 & ~n10432;
  assign n12613 = ~n10429 & n12612;
  assign n12614 = n10434 & ~n12613;
  assign n12615 = ~n10430 & n10432;
  assign n12616 = ~n12614 & ~n12615;
  assign n12617 = ~n6369 & ~n10418;
  assign n12618 = ~n10415 & n12617;
  assign n12619 = n10420 & ~n12618;
  assign n12620 = ~n10416 & n10418;
  assign n12621 = ~n12619 & ~n12620;
  assign n12622 = ~n12616 & n12621;
  assign n12623 = n12616 & ~n12621;
  assign n12624 = ~n12622 & ~n12623;
  assign n12625 = ~n12611 & ~n12624;
  assign n12626 = ~n12610 & ~n12622;
  assign n12627 = ~n12623 & n12626;
  assign n12628 = ~n12607 & n12627;
  assign n12629 = ~n12625 & ~n12628;
  assign n12630 = ~n10392 & ~n10406;
  assign n12631 = ~n10378 & ~n12630;
  assign n12632 = ~n10391 & ~n10405;
  assign n12633 = ~n10402 & n12632;
  assign n12634 = ~n10388 & n12633;
  assign n12635 = ~n12631 & ~n12634;
  assign n12636 = ~n6315 & ~n10396;
  assign n12637 = ~n10393 & n12636;
  assign n12638 = n10398 & ~n12637;
  assign n12639 = ~n10394 & n10396;
  assign n12640 = ~n12638 & ~n12639;
  assign n12641 = ~n6343 & ~n10382;
  assign n12642 = ~n10379 & n12641;
  assign n12643 = n10384 & ~n12642;
  assign n12644 = ~n10380 & n10382;
  assign n12645 = ~n12643 & ~n12644;
  assign n12646 = ~n12640 & n12645;
  assign n12647 = n12640 & ~n12645;
  assign n12648 = ~n12646 & ~n12647;
  assign n12649 = ~n12635 & ~n12648;
  assign n12650 = ~n12634 & ~n12646;
  assign n12651 = ~n12647 & n12650;
  assign n12652 = ~n12631 & n12651;
  assign n12653 = ~n12649 & ~n12652;
  assign n12654 = ~n12629 & n12653;
  assign n12655 = n12629 & ~n12653;
  assign n12656 = ~n12654 & ~n12655;
  assign n12657 = ~n12605 & ~n12656;
  assign n12658 = n12605 & n12656;
  assign n12659 = ~n12657 & ~n12658;
  assign n12660 = ~n10332 & ~n10368;
  assign n12661 = ~n10296 & ~n12660;
  assign n12662 = n10332 & n10368;
  assign n12663 = ~n12661 & ~n12662;
  assign n12664 = ~n10348 & ~n10362;
  assign n12665 = ~n10334 & ~n12664;
  assign n12666 = ~n10347 & ~n10361;
  assign n12667 = ~n10358 & n12666;
  assign n12668 = ~n10344 & n12667;
  assign n12669 = ~n12665 & ~n12668;
  assign n12670 = ~n6451 & ~n10352;
  assign n12671 = ~n10349 & n12670;
  assign n12672 = n10354 & ~n12671;
  assign n12673 = ~n10350 & n10352;
  assign n12674 = ~n12672 & ~n12673;
  assign n12675 = ~n6436 & ~n10338;
  assign n12676 = ~n10335 & n12675;
  assign n12677 = n10340 & ~n12676;
  assign n12678 = ~n10336 & n10338;
  assign n12679 = ~n12677 & ~n12678;
  assign n12680 = ~n12674 & n12679;
  assign n12681 = n12674 & ~n12679;
  assign n12682 = ~n12680 & ~n12681;
  assign n12683 = ~n12669 & ~n12682;
  assign n12684 = ~n12668 & ~n12680;
  assign n12685 = ~n12681 & n12684;
  assign n12686 = ~n12665 & n12685;
  assign n12687 = ~n12683 & ~n12686;
  assign n12688 = ~n10312 & ~n10326;
  assign n12689 = ~n10298 & ~n12688;
  assign n12690 = ~n10311 & ~n10325;
  assign n12691 = ~n10322 & n12690;
  assign n12692 = ~n10308 & n12691;
  assign n12693 = ~n12689 & ~n12692;
  assign n12694 = ~n6487 & ~n10316;
  assign n12695 = ~n10313 & n12694;
  assign n12696 = n10318 & ~n12695;
  assign n12697 = ~n10314 & n10316;
  assign n12698 = ~n12696 & ~n12697;
  assign n12699 = ~n6515 & ~n10302;
  assign n12700 = ~n10299 & n12699;
  assign n12701 = n10304 & ~n12700;
  assign n12702 = ~n10300 & n10302;
  assign n12703 = ~n12701 & ~n12702;
  assign n12704 = ~n12698 & n12703;
  assign n12705 = n12698 & ~n12703;
  assign n12706 = ~n12704 & ~n12705;
  assign n12707 = ~n12693 & ~n12706;
  assign n12708 = ~n12692 & ~n12704;
  assign n12709 = ~n12705 & n12708;
  assign n12710 = ~n12689 & n12709;
  assign n12711 = ~n12707 & ~n12710;
  assign n12712 = ~n12687 & n12711;
  assign n12713 = n12687 & ~n12711;
  assign n12714 = ~n12712 & ~n12713;
  assign n12715 = ~n12663 & ~n12714;
  assign n12716 = n12663 & n12714;
  assign n12717 = ~n12715 & ~n12716;
  assign n12718 = ~n12659 & n12717;
  assign n12719 = n12659 & ~n12717;
  assign n12720 = ~n12718 & ~n12719;
  assign n12721 = ~n12601 & ~n12720;
  assign n12722 = n12601 & n12720;
  assign n12723 = ~n12721 & ~n12722;
  assign n12724 = ~n12597 & n12723;
  assign n12725 = ~n12595 & ~n12723;
  assign n12726 = ~n12596 & n12725;
  assign n12727 = ~n12724 & ~n12726;
  assign n12728 = ~n12414 & ~n12727;
  assign n12729 = n12414 & n12727;
  assign n12730 = ~n12728 & ~n12729;
  assign n12731 = ~n12409 & n12730;
  assign n12732 = n12409 & ~n12730;
  assign n12733 = ~n12731 & ~n12732;
  assign n12734 = ~n11875 & ~n12733;
  assign n12735 = n11875 & n12733;
  assign n12736 = ~n12734 & ~n12735;
  assign n12737 = ~n11516 & ~n11860;
  assign n12738 = ~n11172 & ~n12737;
  assign n12739 = n11516 & n11860;
  assign n12740 = ~n12738 & ~n12739;
  assign n12741 = ~n11686 & ~n11854;
  assign n12742 = ~n11518 & ~n12741;
  assign n12743 = n11686 & n11854;
  assign n12744 = ~n12742 & ~n12743;
  assign n12745 = ~n11768 & ~n11848;
  assign n12746 = ~n11688 & ~n12745;
  assign n12747 = n11768 & n11848;
  assign n12748 = ~n12746 & ~n12747;
  assign n12749 = ~n11806 & ~n11842;
  assign n12750 = ~n11770 & ~n12749;
  assign n12751 = n11806 & n11842;
  assign n12752 = ~n12750 & ~n12751;
  assign n12753 = ~n11822 & ~n11836;
  assign n12754 = ~n11808 & ~n12753;
  assign n12755 = ~n11821 & ~n11835;
  assign n12756 = ~n11832 & n12755;
  assign n12757 = ~n11818 & n12756;
  assign n12758 = ~n12754 & ~n12757;
  assign n12759 = ~n2645 & ~n11826;
  assign n12760 = ~n11823 & n12759;
  assign n12761 = n11828 & ~n12760;
  assign n12762 = ~n11824 & n11826;
  assign n12763 = ~n12761 & ~n12762;
  assign n12764 = ~n2560 & ~n11812;
  assign n12765 = ~n11809 & n12764;
  assign n12766 = n11814 & ~n12765;
  assign n12767 = ~n11810 & n11812;
  assign n12768 = ~n12766 & ~n12767;
  assign n12769 = ~n12763 & n12768;
  assign n12770 = n12763 & ~n12768;
  assign n12771 = ~n12769 & ~n12770;
  assign n12772 = ~n12758 & ~n12771;
  assign n12773 = ~n12757 & ~n12769;
  assign n12774 = ~n12770 & n12773;
  assign n12775 = ~n12754 & n12774;
  assign n12776 = ~n12772 & ~n12775;
  assign n12777 = ~n11786 & ~n11800;
  assign n12778 = ~n11772 & ~n12777;
  assign n12779 = ~n11785 & ~n11799;
  assign n12780 = ~n11796 & n12779;
  assign n12781 = ~n11782 & n12780;
  assign n12782 = ~n12778 & ~n12781;
  assign n12783 = ~n2356 & ~n11790;
  assign n12784 = ~n11787 & n12783;
  assign n12785 = n11792 & ~n12784;
  assign n12786 = ~n11788 & n11790;
  assign n12787 = ~n12785 & ~n12786;
  assign n12788 = ~n2464 & ~n11776;
  assign n12789 = ~n11773 & n12788;
  assign n12790 = n11778 & ~n12789;
  assign n12791 = ~n11774 & n11776;
  assign n12792 = ~n12790 & ~n12791;
  assign n12793 = ~n12787 & n12792;
  assign n12794 = n12787 & ~n12792;
  assign n12795 = ~n12793 & ~n12794;
  assign n12796 = ~n12782 & ~n12795;
  assign n12797 = ~n12781 & ~n12793;
  assign n12798 = ~n12794 & n12797;
  assign n12799 = ~n12778 & n12798;
  assign n12800 = ~n12796 & ~n12799;
  assign n12801 = ~n12776 & n12800;
  assign n12802 = n12776 & ~n12800;
  assign n12803 = ~n12801 & ~n12802;
  assign n12804 = ~n12752 & ~n12803;
  assign n12805 = n12752 & n12803;
  assign n12806 = ~n12804 & ~n12805;
  assign n12807 = ~n11726 & ~n11762;
  assign n12808 = ~n11690 & ~n12807;
  assign n12809 = n11726 & n11762;
  assign n12810 = ~n12808 & ~n12809;
  assign n12811 = ~n11742 & ~n11756;
  assign n12812 = ~n11728 & ~n12811;
  assign n12813 = ~n11741 & ~n11755;
  assign n12814 = ~n11752 & n12813;
  assign n12815 = ~n11738 & n12814;
  assign n12816 = ~n12812 & ~n12815;
  assign n12817 = ~n2027 & ~n11746;
  assign n12818 = ~n11743 & n12817;
  assign n12819 = n11748 & ~n12818;
  assign n12820 = ~n11744 & n11746;
  assign n12821 = ~n12819 & ~n12820;
  assign n12822 = ~n1942 & ~n11732;
  assign n12823 = ~n11729 & n12822;
  assign n12824 = n11734 & ~n12823;
  assign n12825 = ~n11730 & n11732;
  assign n12826 = ~n12824 & ~n12825;
  assign n12827 = ~n12821 & n12826;
  assign n12828 = n12821 & ~n12826;
  assign n12829 = ~n12827 & ~n12828;
  assign n12830 = ~n12816 & ~n12829;
  assign n12831 = ~n12815 & ~n12827;
  assign n12832 = ~n12828 & n12831;
  assign n12833 = ~n12812 & n12832;
  assign n12834 = ~n12830 & ~n12833;
  assign n12835 = ~n11706 & ~n11720;
  assign n12836 = ~n11692 & ~n12835;
  assign n12837 = ~n11705 & ~n11719;
  assign n12838 = ~n11716 & n12837;
  assign n12839 = ~n11702 & n12838;
  assign n12840 = ~n12836 & ~n12839;
  assign n12841 = ~n2229 & ~n11710;
  assign n12842 = ~n11707 & n12841;
  assign n12843 = n11712 & ~n12842;
  assign n12844 = ~n11708 & n11710;
  assign n12845 = ~n12843 & ~n12844;
  assign n12846 = ~n2257 & ~n11696;
  assign n12847 = ~n11693 & n12846;
  assign n12848 = n11698 & ~n12847;
  assign n12849 = ~n11694 & n11696;
  assign n12850 = ~n12848 & ~n12849;
  assign n12851 = ~n12845 & n12850;
  assign n12852 = n12845 & ~n12850;
  assign n12853 = ~n12851 & ~n12852;
  assign n12854 = ~n12840 & ~n12853;
  assign n12855 = ~n12839 & ~n12851;
  assign n12856 = ~n12852 & n12855;
  assign n12857 = ~n12836 & n12856;
  assign n12858 = ~n12854 & ~n12857;
  assign n12859 = ~n12834 & n12858;
  assign n12860 = n12834 & ~n12858;
  assign n12861 = ~n12859 & ~n12860;
  assign n12862 = ~n12810 & ~n12861;
  assign n12863 = n12810 & n12861;
  assign n12864 = ~n12862 & ~n12863;
  assign n12865 = ~n12806 & n12864;
  assign n12866 = n12806 & ~n12864;
  assign n12867 = ~n12865 & ~n12866;
  assign n12868 = ~n12748 & ~n12867;
  assign n12869 = n12748 & n12867;
  assign n12870 = ~n12868 & ~n12869;
  assign n12871 = ~n11600 & ~n11680;
  assign n12872 = ~n11520 & ~n12871;
  assign n12873 = n11600 & n11680;
  assign n12874 = ~n12872 & ~n12873;
  assign n12875 = ~n11638 & ~n11674;
  assign n12876 = ~n11602 & ~n12875;
  assign n12877 = n11638 & n11674;
  assign n12878 = ~n12876 & ~n12877;
  assign n12879 = ~n11654 & ~n11668;
  assign n12880 = ~n11640 & ~n12879;
  assign n12881 = ~n11653 & ~n11667;
  assign n12882 = ~n11664 & n12881;
  assign n12883 = ~n11650 & n12882;
  assign n12884 = ~n12880 & ~n12883;
  assign n12885 = ~n1373 & ~n11658;
  assign n12886 = ~n11655 & n12885;
  assign n12887 = n11660 & ~n12886;
  assign n12888 = ~n11656 & n11658;
  assign n12889 = ~n12887 & ~n12888;
  assign n12890 = ~n1288 & ~n11644;
  assign n12891 = ~n11641 & n12890;
  assign n12892 = n11646 & ~n12891;
  assign n12893 = ~n11642 & n11644;
  assign n12894 = ~n12892 & ~n12893;
  assign n12895 = ~n12889 & n12894;
  assign n12896 = n12889 & ~n12894;
  assign n12897 = ~n12895 & ~n12896;
  assign n12898 = ~n12884 & ~n12897;
  assign n12899 = ~n12883 & ~n12895;
  assign n12900 = ~n12896 & n12899;
  assign n12901 = ~n12880 & n12900;
  assign n12902 = ~n12898 & ~n12901;
  assign n12903 = ~n11618 & ~n11632;
  assign n12904 = ~n11604 & ~n12903;
  assign n12905 = ~n11617 & ~n11631;
  assign n12906 = ~n11628 & n12905;
  assign n12907 = ~n11614 & n12906;
  assign n12908 = ~n12904 & ~n12907;
  assign n12909 = ~n1084 & ~n11622;
  assign n12910 = ~n11619 & n12909;
  assign n12911 = n11624 & ~n12910;
  assign n12912 = ~n11620 & n11622;
  assign n12913 = ~n12911 & ~n12912;
  assign n12914 = ~n1192 & ~n11608;
  assign n12915 = ~n11605 & n12914;
  assign n12916 = n11610 & ~n12915;
  assign n12917 = ~n11606 & n11608;
  assign n12918 = ~n12916 & ~n12917;
  assign n12919 = ~n12913 & n12918;
  assign n12920 = n12913 & ~n12918;
  assign n12921 = ~n12919 & ~n12920;
  assign n12922 = ~n12908 & ~n12921;
  assign n12923 = ~n12907 & ~n12919;
  assign n12924 = ~n12920 & n12923;
  assign n12925 = ~n12904 & n12924;
  assign n12926 = ~n12922 & ~n12925;
  assign n12927 = ~n12902 & n12926;
  assign n12928 = n12902 & ~n12926;
  assign n12929 = ~n12927 & ~n12928;
  assign n12930 = ~n12878 & ~n12929;
  assign n12931 = n12878 & n12929;
  assign n12932 = ~n12930 & ~n12931;
  assign n12933 = ~n11558 & ~n11594;
  assign n12934 = ~n11522 & ~n12933;
  assign n12935 = n11558 & n11594;
  assign n12936 = ~n12934 & ~n12935;
  assign n12937 = ~n11574 & ~n11588;
  assign n12938 = ~n11560 & ~n12937;
  assign n12939 = ~n11573 & ~n11587;
  assign n12940 = ~n11584 & n12939;
  assign n12941 = ~n11570 & n12940;
  assign n12942 = ~n12938 & ~n12941;
  assign n12943 = ~n1768 & ~n11578;
  assign n12944 = ~n11575 & n12943;
  assign n12945 = n11580 & ~n12944;
  assign n12946 = ~n11576 & n11578;
  assign n12947 = ~n12945 & ~n12946;
  assign n12948 = ~n1753 & ~n11564;
  assign n12949 = ~n11561 & n12948;
  assign n12950 = n11566 & ~n12949;
  assign n12951 = ~n11562 & n11564;
  assign n12952 = ~n12950 & ~n12951;
  assign n12953 = ~n12947 & n12952;
  assign n12954 = n12947 & ~n12952;
  assign n12955 = ~n12953 & ~n12954;
  assign n12956 = ~n12942 & ~n12955;
  assign n12957 = ~n12941 & ~n12953;
  assign n12958 = ~n12954 & n12957;
  assign n12959 = ~n12938 & n12958;
  assign n12960 = ~n12956 & ~n12959;
  assign n12961 = ~n11538 & ~n11552;
  assign n12962 = ~n11524 & ~n12961;
  assign n12963 = ~n11537 & ~n11551;
  assign n12964 = ~n11548 & n12963;
  assign n12965 = ~n11534 & n12964;
  assign n12966 = ~n12962 & ~n12965;
  assign n12967 = ~n1804 & ~n11542;
  assign n12968 = ~n11539 & n12967;
  assign n12969 = n11544 & ~n12968;
  assign n12970 = ~n11540 & n11542;
  assign n12971 = ~n12969 & ~n12970;
  assign n12972 = ~n1832 & ~n11528;
  assign n12973 = ~n11525 & n12972;
  assign n12974 = n11530 & ~n12973;
  assign n12975 = ~n11526 & n11528;
  assign n12976 = ~n12974 & ~n12975;
  assign n12977 = ~n12971 & n12976;
  assign n12978 = n12971 & ~n12976;
  assign n12979 = ~n12977 & ~n12978;
  assign n12980 = ~n12966 & ~n12979;
  assign n12981 = ~n12965 & ~n12977;
  assign n12982 = ~n12978 & n12981;
  assign n12983 = ~n12962 & n12982;
  assign n12984 = ~n12980 & ~n12983;
  assign n12985 = ~n12960 & n12984;
  assign n12986 = n12960 & ~n12984;
  assign n12987 = ~n12985 & ~n12986;
  assign n12988 = ~n12936 & ~n12987;
  assign n12989 = n12936 & n12987;
  assign n12990 = ~n12988 & ~n12989;
  assign n12991 = ~n12932 & n12990;
  assign n12992 = n12932 & ~n12990;
  assign n12993 = ~n12991 & ~n12992;
  assign n12994 = ~n12874 & ~n12993;
  assign n12995 = n12874 & n12993;
  assign n12996 = ~n12994 & ~n12995;
  assign n12997 = ~n12870 & n12996;
  assign n12998 = n12870 & ~n12996;
  assign n12999 = ~n12997 & ~n12998;
  assign n13000 = ~n12744 & ~n12999;
  assign n13001 = n12744 & n12999;
  assign n13002 = ~n13000 & ~n13001;
  assign n13003 = ~n11342 & ~n11510;
  assign n13004 = ~n11174 & ~n13003;
  assign n13005 = n11342 & n11510;
  assign n13006 = ~n13004 & ~n13005;
  assign n13007 = ~n11424 & ~n11504;
  assign n13008 = ~n11344 & ~n13007;
  assign n13009 = n11424 & n11504;
  assign n13010 = ~n13008 & ~n13009;
  assign n13011 = ~n11462 & ~n11498;
  assign n13012 = ~n11426 & ~n13011;
  assign n13013 = n11462 & n11498;
  assign n13014 = ~n13012 & ~n13013;
  assign n13015 = ~n11478 & ~n11492;
  assign n13016 = ~n11464 & ~n13015;
  assign n13017 = ~n11477 & ~n11491;
  assign n13018 = ~n11488 & n13017;
  assign n13019 = ~n11474 & n13018;
  assign n13020 = ~n13016 & ~n13019;
  assign n13021 = ~n4174 & ~n11482;
  assign n13022 = ~n11479 & n13021;
  assign n13023 = n11484 & ~n13022;
  assign n13024 = ~n11480 & n11482;
  assign n13025 = ~n13023 & ~n13024;
  assign n13026 = ~n4159 & ~n11468;
  assign n13027 = ~n11465 & n13026;
  assign n13028 = n11470 & ~n13027;
  assign n13029 = ~n11466 & n11468;
  assign n13030 = ~n13028 & ~n13029;
  assign n13031 = ~n13025 & n13030;
  assign n13032 = n13025 & ~n13030;
  assign n13033 = ~n13031 & ~n13032;
  assign n13034 = ~n13020 & ~n13033;
  assign n13035 = ~n13019 & ~n13031;
  assign n13036 = ~n13032 & n13035;
  assign n13037 = ~n13016 & n13036;
  assign n13038 = ~n13034 & ~n13037;
  assign n13039 = ~n11442 & ~n11456;
  assign n13040 = ~n11428 & ~n13039;
  assign n13041 = ~n11441 & ~n11455;
  assign n13042 = ~n11452 & n13041;
  assign n13043 = ~n11438 & n13042;
  assign n13044 = ~n13040 & ~n13043;
  assign n13045 = ~n4105 & ~n11446;
  assign n13046 = ~n11443 & n13045;
  assign n13047 = n11448 & ~n13046;
  assign n13048 = ~n11444 & n11446;
  assign n13049 = ~n13047 & ~n13048;
  assign n13050 = ~n4133 & ~n11432;
  assign n13051 = ~n11429 & n13050;
  assign n13052 = n11434 & ~n13051;
  assign n13053 = ~n11430 & n11432;
  assign n13054 = ~n13052 & ~n13053;
  assign n13055 = ~n13049 & n13054;
  assign n13056 = n13049 & ~n13054;
  assign n13057 = ~n13055 & ~n13056;
  assign n13058 = ~n13044 & ~n13057;
  assign n13059 = ~n13043 & ~n13055;
  assign n13060 = ~n13056 & n13059;
  assign n13061 = ~n13040 & n13060;
  assign n13062 = ~n13058 & ~n13061;
  assign n13063 = ~n13038 & n13062;
  assign n13064 = n13038 & ~n13062;
  assign n13065 = ~n13063 & ~n13064;
  assign n13066 = ~n13014 & ~n13065;
  assign n13067 = n13014 & n13065;
  assign n13068 = ~n13066 & ~n13067;
  assign n13069 = ~n11382 & ~n11418;
  assign n13070 = ~n11346 & ~n13069;
  assign n13071 = n11382 & n11418;
  assign n13072 = ~n13070 & ~n13071;
  assign n13073 = ~n11398 & ~n11412;
  assign n13074 = ~n11384 & ~n13073;
  assign n13075 = ~n11397 & ~n11411;
  assign n13076 = ~n11408 & n13075;
  assign n13077 = ~n11394 & n13076;
  assign n13078 = ~n13074 & ~n13077;
  assign n13079 = ~n4012 & ~n11402;
  assign n13080 = ~n11399 & n13079;
  assign n13081 = n11404 & ~n13080;
  assign n13082 = ~n11400 & n11402;
  assign n13083 = ~n13081 & ~n13082;
  assign n13084 = ~n3997 & ~n11388;
  assign n13085 = ~n11385 & n13084;
  assign n13086 = n11390 & ~n13085;
  assign n13087 = ~n11386 & n11388;
  assign n13088 = ~n13086 & ~n13087;
  assign n13089 = ~n13083 & n13088;
  assign n13090 = n13083 & ~n13088;
  assign n13091 = ~n13089 & ~n13090;
  assign n13092 = ~n13078 & ~n13091;
  assign n13093 = ~n13077 & ~n13089;
  assign n13094 = ~n13090 & n13093;
  assign n13095 = ~n13074 & n13094;
  assign n13096 = ~n13092 & ~n13095;
  assign n13097 = ~n11362 & ~n11376;
  assign n13098 = ~n11348 & ~n13097;
  assign n13099 = ~n11361 & ~n11375;
  assign n13100 = ~n11372 & n13099;
  assign n13101 = ~n11358 & n13100;
  assign n13102 = ~n13098 & ~n13101;
  assign n13103 = ~n4048 & ~n11366;
  assign n13104 = ~n11363 & n13103;
  assign n13105 = n11368 & ~n13104;
  assign n13106 = ~n11364 & n11366;
  assign n13107 = ~n13105 & ~n13106;
  assign n13108 = ~n4076 & ~n11352;
  assign n13109 = ~n11349 & n13108;
  assign n13110 = n11354 & ~n13109;
  assign n13111 = ~n11350 & n11352;
  assign n13112 = ~n13110 & ~n13111;
  assign n13113 = ~n13107 & n13112;
  assign n13114 = n13107 & ~n13112;
  assign n13115 = ~n13113 & ~n13114;
  assign n13116 = ~n13102 & ~n13115;
  assign n13117 = ~n13101 & ~n13113;
  assign n13118 = ~n13114 & n13117;
  assign n13119 = ~n13098 & n13118;
  assign n13120 = ~n13116 & ~n13119;
  assign n13121 = ~n13096 & n13120;
  assign n13122 = n13096 & ~n13120;
  assign n13123 = ~n13121 & ~n13122;
  assign n13124 = ~n13072 & ~n13123;
  assign n13125 = n13072 & n13123;
  assign n13126 = ~n13124 & ~n13125;
  assign n13127 = ~n13068 & n13126;
  assign n13128 = n13068 & ~n13126;
  assign n13129 = ~n13127 & ~n13128;
  assign n13130 = ~n13010 & ~n13129;
  assign n13131 = n13010 & n13129;
  assign n13132 = ~n13130 & ~n13131;
  assign n13133 = ~n11256 & ~n11336;
  assign n13134 = ~n11176 & ~n13133;
  assign n13135 = n11256 & n11336;
  assign n13136 = ~n13134 & ~n13135;
  assign n13137 = ~n11294 & ~n11330;
  assign n13138 = ~n11258 & ~n13137;
  assign n13139 = n11294 & n11330;
  assign n13140 = ~n13138 & ~n13139;
  assign n13141 = ~n11310 & ~n11324;
  assign n13142 = ~n11296 & ~n13141;
  assign n13143 = ~n11309 & ~n11323;
  assign n13144 = ~n11320 & n13143;
  assign n13145 = ~n11306 & n13144;
  assign n13146 = ~n13142 & ~n13145;
  assign n13147 = ~n4303 & ~n11314;
  assign n13148 = ~n11311 & n13147;
  assign n13149 = n11316 & ~n13148;
  assign n13150 = ~n11312 & n11314;
  assign n13151 = ~n13149 & ~n13150;
  assign n13152 = ~n4288 & ~n11300;
  assign n13153 = ~n11297 & n13152;
  assign n13154 = n11302 & ~n13153;
  assign n13155 = ~n11298 & n11300;
  assign n13156 = ~n13154 & ~n13155;
  assign n13157 = ~n13151 & n13156;
  assign n13158 = n13151 & ~n13156;
  assign n13159 = ~n13157 & ~n13158;
  assign n13160 = ~n13146 & ~n13159;
  assign n13161 = ~n13145 & ~n13157;
  assign n13162 = ~n13158 & n13161;
  assign n13163 = ~n13142 & n13162;
  assign n13164 = ~n13160 & ~n13163;
  assign n13165 = ~n11274 & ~n11288;
  assign n13166 = ~n11260 & ~n13165;
  assign n13167 = ~n11273 & ~n11287;
  assign n13168 = ~n11284 & n13167;
  assign n13169 = ~n11270 & n13168;
  assign n13170 = ~n13166 & ~n13169;
  assign n13171 = ~n4234 & ~n11278;
  assign n13172 = ~n11275 & n13171;
  assign n13173 = n11280 & ~n13172;
  assign n13174 = ~n11276 & n11278;
  assign n13175 = ~n13173 & ~n13174;
  assign n13176 = ~n4262 & ~n11264;
  assign n13177 = ~n11261 & n13176;
  assign n13178 = n11266 & ~n13177;
  assign n13179 = ~n11262 & n11264;
  assign n13180 = ~n13178 & ~n13179;
  assign n13181 = ~n13175 & n13180;
  assign n13182 = n13175 & ~n13180;
  assign n13183 = ~n13181 & ~n13182;
  assign n13184 = ~n13170 & ~n13183;
  assign n13185 = ~n13169 & ~n13181;
  assign n13186 = ~n13182 & n13185;
  assign n13187 = ~n13166 & n13186;
  assign n13188 = ~n13184 & ~n13187;
  assign n13189 = ~n13164 & n13188;
  assign n13190 = n13164 & ~n13188;
  assign n13191 = ~n13189 & ~n13190;
  assign n13192 = ~n13140 & ~n13191;
  assign n13193 = n13140 & n13191;
  assign n13194 = ~n13192 & ~n13193;
  assign n13195 = ~n11214 & ~n11250;
  assign n13196 = ~n11178 & ~n13195;
  assign n13197 = n11214 & n11250;
  assign n13198 = ~n13196 & ~n13197;
  assign n13199 = ~n11230 & ~n11244;
  assign n13200 = ~n11216 & ~n13199;
  assign n13201 = ~n11229 & ~n11243;
  assign n13202 = ~n11240 & n13201;
  assign n13203 = ~n11226 & n13202;
  assign n13204 = ~n13200 & ~n13203;
  assign n13205 = ~n4370 & ~n11234;
  assign n13206 = ~n11231 & n13205;
  assign n13207 = n11236 & ~n13206;
  assign n13208 = ~n11232 & n11234;
  assign n13209 = ~n13207 & ~n13208;
  assign n13210 = ~n4355 & ~n11220;
  assign n13211 = ~n11217 & n13210;
  assign n13212 = n11222 & ~n13211;
  assign n13213 = ~n11218 & n11220;
  assign n13214 = ~n13212 & ~n13213;
  assign n13215 = ~n13209 & n13214;
  assign n13216 = n13209 & ~n13214;
  assign n13217 = ~n13215 & ~n13216;
  assign n13218 = ~n13204 & ~n13217;
  assign n13219 = ~n13203 & ~n13215;
  assign n13220 = ~n13216 & n13219;
  assign n13221 = ~n13200 & n13220;
  assign n13222 = ~n13218 & ~n13221;
  assign n13223 = ~n11194 & ~n11208;
  assign n13224 = ~n11180 & ~n13223;
  assign n13225 = ~n11193 & ~n11207;
  assign n13226 = ~n11204 & n13225;
  assign n13227 = ~n11190 & n13226;
  assign n13228 = ~n13224 & ~n13227;
  assign n13229 = ~n4406 & ~n11198;
  assign n13230 = ~n11195 & n13229;
  assign n13231 = n11200 & ~n13230;
  assign n13232 = ~n11196 & n11198;
  assign n13233 = ~n13231 & ~n13232;
  assign n13234 = ~n4434 & ~n11184;
  assign n13235 = ~n11181 & n13234;
  assign n13236 = n11186 & ~n13235;
  assign n13237 = ~n11182 & n11184;
  assign n13238 = ~n13236 & ~n13237;
  assign n13239 = ~n13233 & n13238;
  assign n13240 = n13233 & ~n13238;
  assign n13241 = ~n13239 & ~n13240;
  assign n13242 = ~n13228 & ~n13241;
  assign n13243 = ~n13227 & ~n13239;
  assign n13244 = ~n13240 & n13243;
  assign n13245 = ~n13224 & n13244;
  assign n13246 = ~n13242 & ~n13245;
  assign n13247 = ~n13222 & n13246;
  assign n13248 = n13222 & ~n13246;
  assign n13249 = ~n13247 & ~n13248;
  assign n13250 = ~n13198 & ~n13249;
  assign n13251 = n13198 & n13249;
  assign n13252 = ~n13250 & ~n13251;
  assign n13253 = ~n13194 & n13252;
  assign n13254 = n13194 & ~n13252;
  assign n13255 = ~n13253 & ~n13254;
  assign n13256 = ~n13136 & ~n13255;
  assign n13257 = n13136 & n13255;
  assign n13258 = ~n13256 & ~n13257;
  assign n13259 = ~n13132 & n13258;
  assign n13260 = n13132 & ~n13258;
  assign n13261 = ~n13259 & ~n13260;
  assign n13262 = ~n13006 & ~n13261;
  assign n13263 = n13006 & n13261;
  assign n13264 = ~n13262 & ~n13263;
  assign n13265 = ~n13002 & n13264;
  assign n13266 = n13002 & ~n13264;
  assign n13267 = ~n13265 & ~n13266;
  assign n13268 = ~n12740 & ~n13267;
  assign n13269 = n12740 & n13267;
  assign n13270 = ~n13268 & ~n13269;
  assign n13271 = ~n12736 & ~n13270;
  assign n13272 = ~n11871 & ~n13271;
  assign n13273 = ~n12734 & n13270;
  assign n13274 = ~n12735 & n13273;
  assign n13275 = ~n13272 & ~n13274;
  assign n13276 = ~n12409 & ~n12730;
  assign n13277 = ~n11875 & ~n13276;
  assign n13278 = n12409 & n12730;
  assign n13279 = ~n13277 & ~n13278;
  assign n13280 = ~n12597 & ~n12723;
  assign n13281 = ~n12414 & ~n13280;
  assign n13282 = ~n12595 & n12723;
  assign n13283 = ~n12596 & n13282;
  assign n13284 = ~n13281 & ~n13283;
  assign n13285 = ~n12532 & ~n12590;
  assign n13286 = ~n12419 & ~n13285;
  assign n13287 = ~n12530 & n12590;
  assign n13288 = ~n12531 & n13287;
  assign n13289 = ~n13286 & ~n13288;
  assign n13290 = ~n12481 & ~n12526;
  assign n13291 = ~n12423 & ~n13290;
  assign n13292 = n12481 & n12526;
  assign n13293 = ~n13291 & ~n13292;
  assign n13294 = ~n12486 & ~n12521;
  assign n13295 = ~n12522 & ~n13294;
  assign n13296 = n12507 & n12512;
  assign n13297 = ~n12502 & ~n13296;
  assign n13298 = ~n12507 & ~n12512;
  assign n13299 = ~n12493 & ~n13298;
  assign n13300 = ~n13297 & n13299;
  assign n13301 = ~n13297 & ~n13298;
  assign n13302 = n12493 & ~n13301;
  assign n13303 = ~n13300 & ~n13302;
  assign n13304 = ~n13295 & n13303;
  assign n13305 = ~n12522 & ~n13303;
  assign n13306 = ~n13294 & n13305;
  assign n13307 = ~n13304 & ~n13306;
  assign n13308 = ~n12451 & ~n12475;
  assign n13309 = ~n12427 & ~n13308;
  assign n13310 = ~n12450 & ~n12474;
  assign n13311 = ~n12471 & n13310;
  assign n13312 = ~n12447 & n13311;
  assign n13313 = ~n13309 & ~n13312;
  assign n13314 = n12438 & n12443;
  assign n13315 = ~n12433 & ~n13314;
  assign n13316 = ~n12438 & ~n12443;
  assign n13317 = ~n13315 & ~n13316;
  assign n13318 = n12462 & n12467;
  assign n13319 = ~n12457 & ~n13318;
  assign n13320 = ~n12462 & ~n12467;
  assign n13321 = ~n13319 & ~n13320;
  assign n13322 = ~n13317 & n13321;
  assign n13323 = n13317 & ~n13321;
  assign n13324 = ~n13322 & ~n13323;
  assign n13325 = ~n13313 & ~n13324;
  assign n13326 = ~n13312 & ~n13322;
  assign n13327 = ~n13323 & n13326;
  assign n13328 = ~n13309 & n13327;
  assign n13329 = ~n13325 & ~n13328;
  assign n13330 = ~n13307 & n13329;
  assign n13331 = n13307 & ~n13329;
  assign n13332 = ~n13330 & ~n13331;
  assign n13333 = n13293 & n13332;
  assign n13334 = ~n13293 & ~n13332;
  assign n13335 = ~n12560 & ~n12584;
  assign n13336 = ~n12536 & ~n13335;
  assign n13337 = ~n12559 & ~n12583;
  assign n13338 = ~n12580 & n13337;
  assign n13339 = ~n12556 & n13338;
  assign n13340 = ~n13336 & ~n13339;
  assign n13341 = n12547 & n12552;
  assign n13342 = ~n12542 & ~n13341;
  assign n13343 = ~n12547 & ~n12552;
  assign n13344 = ~n13342 & ~n13343;
  assign n13345 = n12571 & n12576;
  assign n13346 = ~n12566 & ~n13345;
  assign n13347 = ~n12571 & ~n12576;
  assign n13348 = ~n13346 & ~n13347;
  assign n13349 = ~n13344 & n13348;
  assign n13350 = n13344 & ~n13348;
  assign n13351 = ~n13349 & ~n13350;
  assign n13352 = ~n13340 & ~n13351;
  assign n13353 = ~n13339 & ~n13349;
  assign n13354 = ~n13350 & n13353;
  assign n13355 = ~n13336 & n13354;
  assign n13356 = ~n13352 & ~n13355;
  assign n13357 = ~n13334 & ~n13356;
  assign n13358 = ~n13333 & n13357;
  assign n13359 = ~n13333 & ~n13334;
  assign n13360 = n13356 & ~n13359;
  assign n13361 = ~n13358 & ~n13360;
  assign n13362 = n13289 & n13361;
  assign n13363 = ~n13289 & ~n13361;
  assign n13364 = ~n12659 & ~n12717;
  assign n13365 = ~n12601 & ~n13364;
  assign n13366 = n12659 & n12717;
  assign n13367 = ~n13365 & ~n13366;
  assign n13368 = ~n12687 & ~n12711;
  assign n13369 = ~n12663 & ~n13368;
  assign n13370 = ~n12686 & ~n12710;
  assign n13371 = ~n12707 & n13370;
  assign n13372 = ~n12683 & n13371;
  assign n13373 = ~n13369 & ~n13372;
  assign n13374 = n12674 & n12679;
  assign n13375 = ~n12669 & ~n13374;
  assign n13376 = ~n12674 & ~n12679;
  assign n13377 = ~n13375 & ~n13376;
  assign n13378 = n12698 & n12703;
  assign n13379 = ~n12693 & ~n13378;
  assign n13380 = ~n12698 & ~n12703;
  assign n13381 = ~n13379 & ~n13380;
  assign n13382 = ~n13377 & n13381;
  assign n13383 = n13377 & ~n13381;
  assign n13384 = ~n13382 & ~n13383;
  assign n13385 = ~n13373 & ~n13384;
  assign n13386 = ~n13372 & ~n13382;
  assign n13387 = ~n13383 & n13386;
  assign n13388 = ~n13369 & n13387;
  assign n13389 = ~n13385 & ~n13388;
  assign n13390 = ~n12629 & ~n12653;
  assign n13391 = ~n12605 & ~n13390;
  assign n13392 = ~n12628 & ~n12652;
  assign n13393 = ~n12649 & n13392;
  assign n13394 = ~n12625 & n13393;
  assign n13395 = ~n13391 & ~n13394;
  assign n13396 = n12616 & n12621;
  assign n13397 = ~n12611 & ~n13396;
  assign n13398 = ~n12616 & ~n12621;
  assign n13399 = ~n13397 & ~n13398;
  assign n13400 = n12640 & n12645;
  assign n13401 = ~n12635 & ~n13400;
  assign n13402 = ~n12640 & ~n12645;
  assign n13403 = ~n13401 & ~n13402;
  assign n13404 = ~n13399 & n13403;
  assign n13405 = n13399 & ~n13403;
  assign n13406 = ~n13404 & ~n13405;
  assign n13407 = ~n13395 & ~n13406;
  assign n13408 = ~n13394 & ~n13404;
  assign n13409 = ~n13405 & n13408;
  assign n13410 = ~n13391 & n13409;
  assign n13411 = ~n13407 & ~n13410;
  assign n13412 = ~n13389 & n13411;
  assign n13413 = n13389 & ~n13411;
  assign n13414 = ~n13412 & ~n13413;
  assign n13415 = ~n13367 & ~n13414;
  assign n13416 = n13367 & n13414;
  assign n13417 = ~n13415 & ~n13416;
  assign n13418 = ~n13363 & ~n13417;
  assign n13419 = ~n13362 & n13418;
  assign n13420 = ~n13362 & ~n13363;
  assign n13421 = n13417 & ~n13420;
  assign n13422 = ~n13419 & ~n13421;
  assign n13423 = ~n13284 & ~n13422;
  assign n13424 = n13284 & n13422;
  assign n13425 = ~n13423 & ~n13424;
  assign n13426 = ~n12141 & ~n12403;
  assign n13427 = ~n11879 & ~n13426;
  assign n13428 = n12141 & n12403;
  assign n13429 = ~n13427 & ~n13428;
  assign n13430 = ~n12271 & ~n12397;
  assign n13431 = ~n12145 & ~n13430;
  assign n13432 = n12271 & n12397;
  assign n13433 = ~n13431 & ~n13432;
  assign n13434 = ~n12333 & ~n12391;
  assign n13435 = ~n12275 & ~n13434;
  assign n13436 = n12333 & n12391;
  assign n13437 = ~n13435 & ~n13436;
  assign n13438 = ~n12361 & ~n12385;
  assign n13439 = ~n12337 & ~n13438;
  assign n13440 = ~n12360 & ~n12384;
  assign n13441 = ~n12381 & n13440;
  assign n13442 = ~n12357 & n13441;
  assign n13443 = ~n13439 & ~n13442;
  assign n13444 = n12348 & n12353;
  assign n13445 = ~n12343 & ~n13444;
  assign n13446 = ~n12348 & ~n12353;
  assign n13447 = ~n13445 & ~n13446;
  assign n13448 = n12372 & n12377;
  assign n13449 = ~n12367 & ~n13448;
  assign n13450 = ~n12372 & ~n12377;
  assign n13451 = ~n13449 & ~n13450;
  assign n13452 = ~n13447 & n13451;
  assign n13453 = n13447 & ~n13451;
  assign n13454 = ~n13452 & ~n13453;
  assign n13455 = ~n13443 & ~n13454;
  assign n13456 = ~n13442 & ~n13452;
  assign n13457 = ~n13453 & n13456;
  assign n13458 = ~n13439 & n13457;
  assign n13459 = ~n13455 & ~n13458;
  assign n13460 = ~n12303 & ~n12327;
  assign n13461 = ~n12279 & ~n13460;
  assign n13462 = ~n12302 & ~n12326;
  assign n13463 = ~n12323 & n13462;
  assign n13464 = ~n12299 & n13463;
  assign n13465 = ~n13461 & ~n13464;
  assign n13466 = n12290 & n12295;
  assign n13467 = ~n12285 & ~n13466;
  assign n13468 = ~n12290 & ~n12295;
  assign n13469 = ~n13467 & ~n13468;
  assign n13470 = n12314 & n12319;
  assign n13471 = ~n12309 & ~n13470;
  assign n13472 = ~n12314 & ~n12319;
  assign n13473 = ~n13471 & ~n13472;
  assign n13474 = ~n13469 & n13473;
  assign n13475 = n13469 & ~n13473;
  assign n13476 = ~n13474 & ~n13475;
  assign n13477 = ~n13465 & ~n13476;
  assign n13478 = ~n13464 & ~n13474;
  assign n13479 = ~n13475 & n13478;
  assign n13480 = ~n13461 & n13479;
  assign n13481 = ~n13477 & ~n13480;
  assign n13482 = ~n13459 & n13481;
  assign n13483 = n13459 & ~n13481;
  assign n13484 = ~n13482 & ~n13483;
  assign n13485 = ~n13437 & ~n13484;
  assign n13486 = n13437 & n13484;
  assign n13487 = ~n13485 & ~n13486;
  assign n13488 = ~n12207 & ~n12265;
  assign n13489 = ~n12149 & ~n13488;
  assign n13490 = n12207 & n12265;
  assign n13491 = ~n13489 & ~n13490;
  assign n13492 = ~n12235 & ~n12259;
  assign n13493 = ~n12211 & ~n13492;
  assign n13494 = ~n12234 & ~n12258;
  assign n13495 = ~n12255 & n13494;
  assign n13496 = ~n12231 & n13495;
  assign n13497 = ~n13493 & ~n13496;
  assign n13498 = n12222 & n12227;
  assign n13499 = ~n12217 & ~n13498;
  assign n13500 = ~n12222 & ~n12227;
  assign n13501 = ~n13499 & ~n13500;
  assign n13502 = n12246 & n12251;
  assign n13503 = ~n12241 & ~n13502;
  assign n13504 = ~n12246 & ~n12251;
  assign n13505 = ~n13503 & ~n13504;
  assign n13506 = ~n13501 & n13505;
  assign n13507 = n13501 & ~n13505;
  assign n13508 = ~n13506 & ~n13507;
  assign n13509 = ~n13497 & ~n13508;
  assign n13510 = ~n13496 & ~n13506;
  assign n13511 = ~n13507 & n13510;
  assign n13512 = ~n13493 & n13511;
  assign n13513 = ~n13509 & ~n13512;
  assign n13514 = ~n12177 & ~n12201;
  assign n13515 = ~n12153 & ~n13514;
  assign n13516 = ~n12176 & ~n12200;
  assign n13517 = ~n12197 & n13516;
  assign n13518 = ~n12173 & n13517;
  assign n13519 = ~n13515 & ~n13518;
  assign n13520 = n12164 & n12169;
  assign n13521 = ~n12159 & ~n13520;
  assign n13522 = ~n12164 & ~n12169;
  assign n13523 = ~n13521 & ~n13522;
  assign n13524 = n12188 & n12193;
  assign n13525 = ~n12183 & ~n13524;
  assign n13526 = ~n12188 & ~n12193;
  assign n13527 = ~n13525 & ~n13526;
  assign n13528 = ~n13523 & n13527;
  assign n13529 = n13523 & ~n13527;
  assign n13530 = ~n13528 & ~n13529;
  assign n13531 = ~n13519 & ~n13530;
  assign n13532 = ~n13518 & ~n13528;
  assign n13533 = ~n13529 & n13532;
  assign n13534 = ~n13515 & n13533;
  assign n13535 = ~n13531 & ~n13534;
  assign n13536 = ~n13513 & n13535;
  assign n13537 = n13513 & ~n13535;
  assign n13538 = ~n13536 & ~n13537;
  assign n13539 = ~n13491 & ~n13538;
  assign n13540 = n13491 & n13538;
  assign n13541 = ~n13539 & ~n13540;
  assign n13542 = ~n13487 & n13541;
  assign n13543 = n13487 & ~n13541;
  assign n13544 = ~n13542 & ~n13543;
  assign n13545 = ~n13433 & ~n13544;
  assign n13546 = n13433 & n13544;
  assign n13547 = ~n13545 & ~n13546;
  assign n13548 = ~n12009 & ~n12135;
  assign n13549 = ~n11883 & ~n13548;
  assign n13550 = n12009 & n12135;
  assign n13551 = ~n13549 & ~n13550;
  assign n13552 = ~n12071 & ~n12129;
  assign n13553 = ~n12013 & ~n13552;
  assign n13554 = n12071 & n12129;
  assign n13555 = ~n13553 & ~n13554;
  assign n13556 = ~n12099 & ~n12123;
  assign n13557 = ~n12075 & ~n13556;
  assign n13558 = ~n12098 & ~n12122;
  assign n13559 = ~n12119 & n13558;
  assign n13560 = ~n12095 & n13559;
  assign n13561 = ~n13557 & ~n13560;
  assign n13562 = n12086 & n12091;
  assign n13563 = ~n12081 & ~n13562;
  assign n13564 = ~n12086 & ~n12091;
  assign n13565 = ~n13563 & ~n13564;
  assign n13566 = n12110 & n12115;
  assign n13567 = ~n12105 & ~n13566;
  assign n13568 = ~n12110 & ~n12115;
  assign n13569 = ~n13567 & ~n13568;
  assign n13570 = ~n13565 & n13569;
  assign n13571 = n13565 & ~n13569;
  assign n13572 = ~n13570 & ~n13571;
  assign n13573 = ~n13561 & ~n13572;
  assign n13574 = ~n13560 & ~n13570;
  assign n13575 = ~n13571 & n13574;
  assign n13576 = ~n13557 & n13575;
  assign n13577 = ~n13573 & ~n13576;
  assign n13578 = ~n12041 & ~n12065;
  assign n13579 = ~n12017 & ~n13578;
  assign n13580 = ~n12040 & ~n12064;
  assign n13581 = ~n12061 & n13580;
  assign n13582 = ~n12037 & n13581;
  assign n13583 = ~n13579 & ~n13582;
  assign n13584 = n12028 & n12033;
  assign n13585 = ~n12023 & ~n13584;
  assign n13586 = ~n12028 & ~n12033;
  assign n13587 = ~n13585 & ~n13586;
  assign n13588 = n12052 & n12057;
  assign n13589 = ~n12047 & ~n13588;
  assign n13590 = ~n12052 & ~n12057;
  assign n13591 = ~n13589 & ~n13590;
  assign n13592 = ~n13587 & n13591;
  assign n13593 = n13587 & ~n13591;
  assign n13594 = ~n13592 & ~n13593;
  assign n13595 = ~n13583 & ~n13594;
  assign n13596 = ~n13582 & ~n13592;
  assign n13597 = ~n13593 & n13596;
  assign n13598 = ~n13579 & n13597;
  assign n13599 = ~n13595 & ~n13598;
  assign n13600 = ~n13577 & n13599;
  assign n13601 = n13577 & ~n13599;
  assign n13602 = ~n13600 & ~n13601;
  assign n13603 = ~n13555 & ~n13602;
  assign n13604 = n13555 & n13602;
  assign n13605 = ~n13603 & ~n13604;
  assign n13606 = ~n11945 & ~n12003;
  assign n13607 = ~n11887 & ~n13606;
  assign n13608 = n11945 & n12003;
  assign n13609 = ~n13607 & ~n13608;
  assign n13610 = ~n11973 & ~n11997;
  assign n13611 = ~n11949 & ~n13610;
  assign n13612 = ~n11972 & ~n11996;
  assign n13613 = ~n11993 & n13612;
  assign n13614 = ~n11969 & n13613;
  assign n13615 = ~n13611 & ~n13614;
  assign n13616 = n11960 & n11965;
  assign n13617 = ~n11955 & ~n13616;
  assign n13618 = ~n11960 & ~n11965;
  assign n13619 = ~n13617 & ~n13618;
  assign n13620 = n11984 & n11989;
  assign n13621 = ~n11979 & ~n13620;
  assign n13622 = ~n11984 & ~n11989;
  assign n13623 = ~n13621 & ~n13622;
  assign n13624 = ~n13619 & n13623;
  assign n13625 = n13619 & ~n13623;
  assign n13626 = ~n13624 & ~n13625;
  assign n13627 = ~n13615 & ~n13626;
  assign n13628 = ~n13614 & ~n13624;
  assign n13629 = ~n13625 & n13628;
  assign n13630 = ~n13611 & n13629;
  assign n13631 = ~n13627 & ~n13630;
  assign n13632 = ~n11915 & ~n11939;
  assign n13633 = ~n11891 & ~n13632;
  assign n13634 = ~n11914 & ~n11938;
  assign n13635 = ~n11935 & n13634;
  assign n13636 = ~n11911 & n13635;
  assign n13637 = ~n13633 & ~n13636;
  assign n13638 = n11902 & n11907;
  assign n13639 = ~n11897 & ~n13638;
  assign n13640 = ~n11902 & ~n11907;
  assign n13641 = ~n13639 & ~n13640;
  assign n13642 = n11926 & n11931;
  assign n13643 = ~n11921 & ~n13642;
  assign n13644 = ~n11926 & ~n11931;
  assign n13645 = ~n13643 & ~n13644;
  assign n13646 = ~n13641 & n13645;
  assign n13647 = n13641 & ~n13645;
  assign n13648 = ~n13646 & ~n13647;
  assign n13649 = ~n13637 & ~n13648;
  assign n13650 = ~n13636 & ~n13646;
  assign n13651 = ~n13647 & n13650;
  assign n13652 = ~n13633 & n13651;
  assign n13653 = ~n13649 & ~n13652;
  assign n13654 = ~n13631 & n13653;
  assign n13655 = n13631 & ~n13653;
  assign n13656 = ~n13654 & ~n13655;
  assign n13657 = ~n13609 & ~n13656;
  assign n13658 = n13609 & n13656;
  assign n13659 = ~n13657 & ~n13658;
  assign n13660 = ~n13605 & n13659;
  assign n13661 = n13605 & ~n13659;
  assign n13662 = ~n13660 & ~n13661;
  assign n13663 = ~n13551 & ~n13662;
  assign n13664 = n13551 & n13662;
  assign n13665 = ~n13663 & ~n13664;
  assign n13666 = ~n13547 & n13665;
  assign n13667 = n13547 & ~n13665;
  assign n13668 = ~n13666 & ~n13667;
  assign n13669 = ~n13429 & ~n13668;
  assign n13670 = n13429 & n13668;
  assign n13671 = ~n13669 & ~n13670;
  assign n13672 = ~n13425 & n13671;
  assign n13673 = n13425 & ~n13671;
  assign n13674 = ~n13672 & ~n13673;
  assign n13675 = ~n13279 & ~n13674;
  assign n13676 = n13279 & n13674;
  assign n13677 = ~n13675 & ~n13676;
  assign n13678 = ~n13002 & ~n13264;
  assign n13679 = ~n12740 & ~n13678;
  assign n13680 = n13002 & n13264;
  assign n13681 = ~n13679 & ~n13680;
  assign n13682 = ~n13132 & ~n13258;
  assign n13683 = ~n13006 & ~n13682;
  assign n13684 = n13132 & n13258;
  assign n13685 = ~n13683 & ~n13684;
  assign n13686 = ~n13194 & ~n13252;
  assign n13687 = ~n13136 & ~n13686;
  assign n13688 = n13194 & n13252;
  assign n13689 = ~n13687 & ~n13688;
  assign n13690 = ~n13222 & ~n13246;
  assign n13691 = ~n13198 & ~n13690;
  assign n13692 = ~n13221 & ~n13245;
  assign n13693 = ~n13242 & n13692;
  assign n13694 = ~n13218 & n13693;
  assign n13695 = ~n13691 & ~n13694;
  assign n13696 = n13209 & n13214;
  assign n13697 = ~n13204 & ~n13696;
  assign n13698 = ~n13209 & ~n13214;
  assign n13699 = ~n13697 & ~n13698;
  assign n13700 = n13233 & n13238;
  assign n13701 = ~n13228 & ~n13700;
  assign n13702 = ~n13233 & ~n13238;
  assign n13703 = ~n13701 & ~n13702;
  assign n13704 = ~n13699 & n13703;
  assign n13705 = n13699 & ~n13703;
  assign n13706 = ~n13704 & ~n13705;
  assign n13707 = ~n13695 & ~n13706;
  assign n13708 = ~n13694 & ~n13704;
  assign n13709 = ~n13705 & n13708;
  assign n13710 = ~n13691 & n13709;
  assign n13711 = ~n13707 & ~n13710;
  assign n13712 = ~n13164 & ~n13188;
  assign n13713 = ~n13140 & ~n13712;
  assign n13714 = ~n13163 & ~n13187;
  assign n13715 = ~n13184 & n13714;
  assign n13716 = ~n13160 & n13715;
  assign n13717 = ~n13713 & ~n13716;
  assign n13718 = n13151 & n13156;
  assign n13719 = ~n13146 & ~n13718;
  assign n13720 = ~n13151 & ~n13156;
  assign n13721 = ~n13719 & ~n13720;
  assign n13722 = n13175 & n13180;
  assign n13723 = ~n13170 & ~n13722;
  assign n13724 = ~n13175 & ~n13180;
  assign n13725 = ~n13723 & ~n13724;
  assign n13726 = ~n13721 & n13725;
  assign n13727 = n13721 & ~n13725;
  assign n13728 = ~n13726 & ~n13727;
  assign n13729 = ~n13717 & ~n13728;
  assign n13730 = ~n13716 & ~n13726;
  assign n13731 = ~n13727 & n13730;
  assign n13732 = ~n13713 & n13731;
  assign n13733 = ~n13729 & ~n13732;
  assign n13734 = ~n13711 & n13733;
  assign n13735 = n13711 & ~n13733;
  assign n13736 = ~n13734 & ~n13735;
  assign n13737 = ~n13689 & ~n13736;
  assign n13738 = n13689 & n13736;
  assign n13739 = ~n13737 & ~n13738;
  assign n13740 = ~n13068 & ~n13126;
  assign n13741 = ~n13010 & ~n13740;
  assign n13742 = n13068 & n13126;
  assign n13743 = ~n13741 & ~n13742;
  assign n13744 = ~n13096 & ~n13120;
  assign n13745 = ~n13072 & ~n13744;
  assign n13746 = ~n13095 & ~n13119;
  assign n13747 = ~n13116 & n13746;
  assign n13748 = ~n13092 & n13747;
  assign n13749 = ~n13745 & ~n13748;
  assign n13750 = n13083 & n13088;
  assign n13751 = ~n13078 & ~n13750;
  assign n13752 = ~n13083 & ~n13088;
  assign n13753 = ~n13751 & ~n13752;
  assign n13754 = n13107 & n13112;
  assign n13755 = ~n13102 & ~n13754;
  assign n13756 = ~n13107 & ~n13112;
  assign n13757 = ~n13755 & ~n13756;
  assign n13758 = ~n13753 & n13757;
  assign n13759 = n13753 & ~n13757;
  assign n13760 = ~n13758 & ~n13759;
  assign n13761 = ~n13749 & ~n13760;
  assign n13762 = ~n13748 & ~n13758;
  assign n13763 = ~n13759 & n13762;
  assign n13764 = ~n13745 & n13763;
  assign n13765 = ~n13761 & ~n13764;
  assign n13766 = ~n13038 & ~n13062;
  assign n13767 = ~n13014 & ~n13766;
  assign n13768 = ~n13037 & ~n13061;
  assign n13769 = ~n13058 & n13768;
  assign n13770 = ~n13034 & n13769;
  assign n13771 = ~n13767 & ~n13770;
  assign n13772 = n13025 & n13030;
  assign n13773 = ~n13020 & ~n13772;
  assign n13774 = ~n13025 & ~n13030;
  assign n13775 = ~n13773 & ~n13774;
  assign n13776 = n13049 & n13054;
  assign n13777 = ~n13044 & ~n13776;
  assign n13778 = ~n13049 & ~n13054;
  assign n13779 = ~n13777 & ~n13778;
  assign n13780 = ~n13775 & n13779;
  assign n13781 = n13775 & ~n13779;
  assign n13782 = ~n13780 & ~n13781;
  assign n13783 = ~n13771 & ~n13782;
  assign n13784 = ~n13770 & ~n13780;
  assign n13785 = ~n13781 & n13784;
  assign n13786 = ~n13767 & n13785;
  assign n13787 = ~n13783 & ~n13786;
  assign n13788 = ~n13765 & n13787;
  assign n13789 = n13765 & ~n13787;
  assign n13790 = ~n13788 & ~n13789;
  assign n13791 = ~n13743 & ~n13790;
  assign n13792 = n13743 & n13790;
  assign n13793 = ~n13791 & ~n13792;
  assign n13794 = ~n13739 & n13793;
  assign n13795 = n13739 & ~n13793;
  assign n13796 = ~n13794 & ~n13795;
  assign n13797 = ~n13685 & ~n13796;
  assign n13798 = n13685 & n13796;
  assign n13799 = ~n13797 & ~n13798;
  assign n13800 = ~n12870 & ~n12996;
  assign n13801 = ~n12744 & ~n13800;
  assign n13802 = n12870 & n12996;
  assign n13803 = ~n13801 & ~n13802;
  assign n13804 = ~n12932 & ~n12990;
  assign n13805 = ~n12874 & ~n13804;
  assign n13806 = n12932 & n12990;
  assign n13807 = ~n13805 & ~n13806;
  assign n13808 = ~n12960 & ~n12984;
  assign n13809 = ~n12936 & ~n13808;
  assign n13810 = ~n12959 & ~n12983;
  assign n13811 = ~n12980 & n13810;
  assign n13812 = ~n12956 & n13811;
  assign n13813 = ~n13809 & ~n13812;
  assign n13814 = n12947 & n12952;
  assign n13815 = ~n12942 & ~n13814;
  assign n13816 = ~n12947 & ~n12952;
  assign n13817 = ~n13815 & ~n13816;
  assign n13818 = n12971 & n12976;
  assign n13819 = ~n12966 & ~n13818;
  assign n13820 = ~n12971 & ~n12976;
  assign n13821 = ~n13819 & ~n13820;
  assign n13822 = ~n13817 & n13821;
  assign n13823 = n13817 & ~n13821;
  assign n13824 = ~n13822 & ~n13823;
  assign n13825 = ~n13813 & ~n13824;
  assign n13826 = ~n13812 & ~n13822;
  assign n13827 = ~n13823 & n13826;
  assign n13828 = ~n13809 & n13827;
  assign n13829 = ~n13825 & ~n13828;
  assign n13830 = ~n12902 & ~n12926;
  assign n13831 = ~n12878 & ~n13830;
  assign n13832 = ~n12901 & ~n12925;
  assign n13833 = ~n12922 & n13832;
  assign n13834 = ~n12898 & n13833;
  assign n13835 = ~n13831 & ~n13834;
  assign n13836 = n12889 & n12894;
  assign n13837 = ~n12884 & ~n13836;
  assign n13838 = ~n12889 & ~n12894;
  assign n13839 = ~n13837 & ~n13838;
  assign n13840 = n12913 & n12918;
  assign n13841 = ~n12908 & ~n13840;
  assign n13842 = ~n12913 & ~n12918;
  assign n13843 = ~n13841 & ~n13842;
  assign n13844 = ~n13839 & n13843;
  assign n13845 = n13839 & ~n13843;
  assign n13846 = ~n13844 & ~n13845;
  assign n13847 = ~n13835 & ~n13846;
  assign n13848 = ~n13834 & ~n13844;
  assign n13849 = ~n13845 & n13848;
  assign n13850 = ~n13831 & n13849;
  assign n13851 = ~n13847 & ~n13850;
  assign n13852 = ~n13829 & n13851;
  assign n13853 = n13829 & ~n13851;
  assign n13854 = ~n13852 & ~n13853;
  assign n13855 = ~n13807 & ~n13854;
  assign n13856 = n13807 & n13854;
  assign n13857 = ~n13855 & ~n13856;
  assign n13858 = ~n12806 & ~n12864;
  assign n13859 = ~n12748 & ~n13858;
  assign n13860 = n12806 & n12864;
  assign n13861 = ~n13859 & ~n13860;
  assign n13862 = ~n12834 & ~n12858;
  assign n13863 = ~n12810 & ~n13862;
  assign n13864 = ~n12833 & ~n12857;
  assign n13865 = ~n12854 & n13864;
  assign n13866 = ~n12830 & n13865;
  assign n13867 = ~n13863 & ~n13866;
  assign n13868 = n12821 & n12826;
  assign n13869 = ~n12816 & ~n13868;
  assign n13870 = ~n12821 & ~n12826;
  assign n13871 = ~n13869 & ~n13870;
  assign n13872 = n12845 & n12850;
  assign n13873 = ~n12840 & ~n13872;
  assign n13874 = ~n12845 & ~n12850;
  assign n13875 = ~n13873 & ~n13874;
  assign n13876 = ~n13871 & n13875;
  assign n13877 = n13871 & ~n13875;
  assign n13878 = ~n13876 & ~n13877;
  assign n13879 = ~n13867 & ~n13878;
  assign n13880 = ~n13866 & ~n13876;
  assign n13881 = ~n13877 & n13880;
  assign n13882 = ~n13863 & n13881;
  assign n13883 = ~n13879 & ~n13882;
  assign n13884 = ~n12776 & ~n12800;
  assign n13885 = ~n12752 & ~n13884;
  assign n13886 = ~n12775 & ~n12799;
  assign n13887 = ~n12796 & n13886;
  assign n13888 = ~n12772 & n13887;
  assign n13889 = ~n13885 & ~n13888;
  assign n13890 = n12763 & n12768;
  assign n13891 = ~n12758 & ~n13890;
  assign n13892 = ~n12763 & ~n12768;
  assign n13893 = ~n13891 & ~n13892;
  assign n13894 = n12787 & n12792;
  assign n13895 = ~n12782 & ~n13894;
  assign n13896 = ~n12787 & ~n12792;
  assign n13897 = ~n13895 & ~n13896;
  assign n13898 = ~n13893 & n13897;
  assign n13899 = n13893 & ~n13897;
  assign n13900 = ~n13898 & ~n13899;
  assign n13901 = ~n13889 & ~n13900;
  assign n13902 = ~n13888 & ~n13898;
  assign n13903 = ~n13899 & n13902;
  assign n13904 = ~n13885 & n13903;
  assign n13905 = ~n13901 & ~n13904;
  assign n13906 = ~n13883 & n13905;
  assign n13907 = n13883 & ~n13905;
  assign n13908 = ~n13906 & ~n13907;
  assign n13909 = ~n13861 & ~n13908;
  assign n13910 = n13861 & n13908;
  assign n13911 = ~n13909 & ~n13910;
  assign n13912 = ~n13857 & n13911;
  assign n13913 = n13857 & ~n13911;
  assign n13914 = ~n13912 & ~n13913;
  assign n13915 = ~n13803 & ~n13914;
  assign n13916 = n13803 & n13914;
  assign n13917 = ~n13915 & ~n13916;
  assign n13918 = ~n13799 & n13917;
  assign n13919 = n13799 & ~n13917;
  assign n13920 = ~n13918 & ~n13919;
  assign n13921 = ~n13681 & ~n13920;
  assign n13922 = n13681 & n13920;
  assign n13923 = ~n13921 & ~n13922;
  assign n13924 = ~n13677 & ~n13923;
  assign n13925 = ~n13275 & ~n13924;
  assign n13926 = ~n13675 & n13923;
  assign n13927 = ~n13676 & n13926;
  assign n13928 = ~n13925 & ~n13927;
  assign n13929 = ~n13425 & ~n13671;
  assign n13930 = ~n13279 & ~n13929;
  assign n13931 = n13425 & n13671;
  assign n13932 = ~n13930 & ~n13931;
  assign n13933 = ~n13547 & ~n13665;
  assign n13934 = ~n13429 & ~n13933;
  assign n13935 = n13547 & n13665;
  assign n13936 = ~n13934 & ~n13935;
  assign n13937 = ~n13605 & ~n13659;
  assign n13938 = ~n13551 & ~n13937;
  assign n13939 = n13605 & n13659;
  assign n13940 = ~n13938 & ~n13939;
  assign n13941 = ~n13631 & ~n13653;
  assign n13942 = ~n13609 & ~n13941;
  assign n13943 = ~n13630 & ~n13652;
  assign n13944 = ~n13649 & n13943;
  assign n13945 = ~n13627 & n13944;
  assign n13946 = ~n13942 & ~n13945;
  assign n13947 = ~n13640 & ~n13644;
  assign n13948 = ~n13643 & n13947;
  assign n13949 = ~n13639 & n13948;
  assign n13950 = ~n13637 & ~n13949;
  assign n13951 = ~n13641 & ~n13645;
  assign n13952 = ~n13950 & ~n13951;
  assign n13953 = ~n13618 & ~n13622;
  assign n13954 = ~n13621 & n13953;
  assign n13955 = ~n13617 & n13954;
  assign n13956 = ~n13615 & ~n13955;
  assign n13957 = ~n13619 & ~n13623;
  assign n13958 = ~n13956 & ~n13957;
  assign n13959 = ~n13952 & n13958;
  assign n13960 = n13952 & ~n13958;
  assign n13961 = ~n13959 & ~n13960;
  assign n13962 = ~n13946 & ~n13961;
  assign n13963 = ~n13945 & ~n13959;
  assign n13964 = ~n13960 & n13963;
  assign n13965 = ~n13942 & n13964;
  assign n13966 = ~n13962 & ~n13965;
  assign n13967 = ~n13577 & ~n13599;
  assign n13968 = ~n13555 & ~n13967;
  assign n13969 = ~n13576 & ~n13598;
  assign n13970 = ~n13595 & n13969;
  assign n13971 = ~n13573 & n13970;
  assign n13972 = ~n13968 & ~n13971;
  assign n13973 = ~n13586 & ~n13590;
  assign n13974 = ~n13589 & n13973;
  assign n13975 = ~n13585 & n13974;
  assign n13976 = ~n13583 & ~n13975;
  assign n13977 = ~n13587 & ~n13591;
  assign n13978 = ~n13976 & ~n13977;
  assign n13979 = ~n13564 & ~n13568;
  assign n13980 = ~n13567 & n13979;
  assign n13981 = ~n13563 & n13980;
  assign n13982 = ~n13561 & ~n13981;
  assign n13983 = ~n13565 & ~n13569;
  assign n13984 = ~n13982 & ~n13983;
  assign n13985 = ~n13978 & n13984;
  assign n13986 = n13978 & ~n13984;
  assign n13987 = ~n13985 & ~n13986;
  assign n13988 = ~n13972 & ~n13987;
  assign n13989 = ~n13971 & ~n13985;
  assign n13990 = ~n13986 & n13989;
  assign n13991 = ~n13968 & n13990;
  assign n13992 = ~n13988 & ~n13991;
  assign n13993 = ~n13966 & n13992;
  assign n13994 = n13966 & ~n13992;
  assign n13995 = ~n13993 & ~n13994;
  assign n13996 = ~n13940 & ~n13995;
  assign n13997 = n13940 & n13995;
  assign n13998 = ~n13996 & ~n13997;
  assign n13999 = ~n13487 & ~n13541;
  assign n14000 = ~n13433 & ~n13999;
  assign n14001 = n13487 & n13541;
  assign n14002 = ~n14000 & ~n14001;
  assign n14003 = ~n13513 & ~n13535;
  assign n14004 = ~n13491 & ~n14003;
  assign n14005 = ~n13512 & ~n13534;
  assign n14006 = ~n13531 & n14005;
  assign n14007 = ~n13509 & n14006;
  assign n14008 = ~n14004 & ~n14007;
  assign n14009 = ~n13522 & ~n13526;
  assign n14010 = ~n13525 & n14009;
  assign n14011 = ~n13521 & n14010;
  assign n14012 = ~n13519 & ~n14011;
  assign n14013 = ~n13523 & ~n13527;
  assign n14014 = ~n14012 & ~n14013;
  assign n14015 = ~n13500 & ~n13504;
  assign n14016 = ~n13503 & n14015;
  assign n14017 = ~n13499 & n14016;
  assign n14018 = ~n13497 & ~n14017;
  assign n14019 = ~n13501 & ~n13505;
  assign n14020 = ~n14018 & ~n14019;
  assign n14021 = ~n14014 & n14020;
  assign n14022 = n14014 & ~n14020;
  assign n14023 = ~n14021 & ~n14022;
  assign n14024 = ~n14008 & ~n14023;
  assign n14025 = ~n14007 & ~n14021;
  assign n14026 = ~n14022 & n14025;
  assign n14027 = ~n14004 & n14026;
  assign n14028 = ~n14024 & ~n14027;
  assign n14029 = ~n13459 & ~n13481;
  assign n14030 = ~n13437 & ~n14029;
  assign n14031 = ~n13458 & ~n13480;
  assign n14032 = ~n13477 & n14031;
  assign n14033 = ~n13455 & n14032;
  assign n14034 = ~n14030 & ~n14033;
  assign n14035 = ~n13468 & ~n13472;
  assign n14036 = ~n13471 & n14035;
  assign n14037 = ~n13467 & n14036;
  assign n14038 = ~n13465 & ~n14037;
  assign n14039 = ~n13469 & ~n13473;
  assign n14040 = ~n14038 & ~n14039;
  assign n14041 = ~n13446 & ~n13450;
  assign n14042 = ~n13449 & n14041;
  assign n14043 = ~n13445 & n14042;
  assign n14044 = ~n13443 & ~n14043;
  assign n14045 = ~n13447 & ~n13451;
  assign n14046 = ~n14044 & ~n14045;
  assign n14047 = ~n14040 & n14046;
  assign n14048 = n14040 & ~n14046;
  assign n14049 = ~n14047 & ~n14048;
  assign n14050 = ~n14034 & ~n14049;
  assign n14051 = ~n14033 & ~n14047;
  assign n14052 = ~n14048 & n14051;
  assign n14053 = ~n14030 & n14052;
  assign n14054 = ~n14050 & ~n14053;
  assign n14055 = ~n14028 & n14054;
  assign n14056 = n14028 & ~n14054;
  assign n14057 = ~n14055 & ~n14056;
  assign n14058 = ~n14002 & ~n14057;
  assign n14059 = n14002 & n14057;
  assign n14060 = ~n14058 & ~n14059;
  assign n14061 = ~n13998 & n14060;
  assign n14062 = n13998 & ~n14060;
  assign n14063 = ~n14061 & ~n14062;
  assign n14064 = ~n13936 & ~n14063;
  assign n14065 = n13936 & n14063;
  assign n14066 = ~n14064 & ~n14065;
  assign n14067 = ~n13417 & ~n13420;
  assign n14068 = ~n13284 & ~n14067;
  assign n14069 = ~n13363 & n13417;
  assign n14070 = ~n13362 & n14069;
  assign n14071 = ~n14068 & ~n14070;
  assign n14072 = ~n13356 & ~n13359;
  assign n14073 = ~n13289 & ~n14072;
  assign n14074 = ~n13334 & n13356;
  assign n14075 = ~n13333 & n14074;
  assign n14076 = ~n14073 & ~n14075;
  assign n14077 = ~n13307 & ~n13329;
  assign n14078 = ~n13293 & ~n14077;
  assign n14079 = ~n13306 & ~n13328;
  assign n14080 = ~n13325 & n14079;
  assign n14081 = ~n13304 & n14080;
  assign n14082 = ~n14078 & ~n14081;
  assign n14083 = ~n13316 & ~n13320;
  assign n14084 = ~n13319 & n14083;
  assign n14085 = ~n13315 & n14084;
  assign n14086 = ~n13313 & ~n14085;
  assign n14087 = ~n13317 & ~n13321;
  assign n14088 = ~n14086 & ~n14087;
  assign n14089 = ~n13295 & ~n13300;
  assign n14090 = ~n13302 & ~n14089;
  assign n14091 = ~n14088 & n14090;
  assign n14092 = n14088 & ~n14090;
  assign n14093 = ~n14091 & ~n14092;
  assign n14094 = ~n14082 & ~n14093;
  assign n14095 = ~n14081 & ~n14091;
  assign n14096 = ~n14092 & n14095;
  assign n14097 = ~n14078 & n14096;
  assign n14098 = ~n13343 & ~n13347;
  assign n14099 = ~n13346 & n14098;
  assign n14100 = ~n13342 & n14099;
  assign n14101 = ~n13340 & ~n14100;
  assign n14102 = ~n13344 & ~n13348;
  assign n14103 = ~n14101 & ~n14102;
  assign n14104 = ~n14097 & n14103;
  assign n14105 = ~n14094 & n14104;
  assign n14106 = ~n14094 & ~n14097;
  assign n14107 = ~n14103 & ~n14106;
  assign n14108 = ~n14105 & ~n14107;
  assign n14109 = ~n14076 & ~n14108;
  assign n14110 = ~n14075 & ~n14105;
  assign n14111 = ~n14073 & n14110;
  assign n14112 = ~n14107 & n14111;
  assign n14113 = ~n14109 & ~n14112;
  assign n14114 = ~n13389 & ~n13411;
  assign n14115 = ~n13367 & ~n14114;
  assign n14116 = ~n13388 & ~n13410;
  assign n14117 = ~n13407 & n14116;
  assign n14118 = ~n13385 & n14117;
  assign n14119 = ~n14115 & ~n14118;
  assign n14120 = ~n13398 & ~n13402;
  assign n14121 = ~n13401 & n14120;
  assign n14122 = ~n13397 & n14121;
  assign n14123 = ~n13395 & ~n14122;
  assign n14124 = ~n13399 & ~n13403;
  assign n14125 = ~n14123 & ~n14124;
  assign n14126 = ~n13376 & ~n13380;
  assign n14127 = ~n13379 & n14126;
  assign n14128 = ~n13375 & n14127;
  assign n14129 = ~n13373 & ~n14128;
  assign n14130 = ~n13377 & ~n13381;
  assign n14131 = ~n14129 & ~n14130;
  assign n14132 = ~n14125 & n14131;
  assign n14133 = n14125 & ~n14131;
  assign n14134 = ~n14132 & ~n14133;
  assign n14135 = ~n14119 & ~n14134;
  assign n14136 = ~n14118 & ~n14132;
  assign n14137 = ~n14133 & n14136;
  assign n14138 = ~n14115 & n14137;
  assign n14139 = ~n14135 & ~n14138;
  assign n14140 = ~n14113 & n14139;
  assign n14141 = ~n14109 & ~n14139;
  assign n14142 = ~n14112 & n14141;
  assign n14143 = ~n14140 & ~n14142;
  assign n14144 = ~n14071 & ~n14143;
  assign n14145 = n14071 & n14143;
  assign n14146 = ~n14144 & ~n14145;
  assign n14147 = ~n14066 & n14146;
  assign n14148 = n14066 & ~n14146;
  assign n14149 = ~n14147 & ~n14148;
  assign n14150 = ~n13932 & ~n14149;
  assign n14151 = n13932 & n14149;
  assign n14152 = ~n14150 & ~n14151;
  assign n14153 = ~n13799 & ~n13917;
  assign n14154 = ~n13681 & ~n14153;
  assign n14155 = n13799 & n13917;
  assign n14156 = ~n14154 & ~n14155;
  assign n14157 = ~n13857 & ~n13911;
  assign n14158 = ~n13803 & ~n14157;
  assign n14159 = n13857 & n13911;
  assign n14160 = ~n14158 & ~n14159;
  assign n14161 = ~n13883 & ~n13905;
  assign n14162 = ~n13861 & ~n14161;
  assign n14163 = ~n13882 & ~n13904;
  assign n14164 = ~n13901 & n14163;
  assign n14165 = ~n13879 & n14164;
  assign n14166 = ~n14162 & ~n14165;
  assign n14167 = ~n13892 & ~n13896;
  assign n14168 = ~n13895 & n14167;
  assign n14169 = ~n13891 & n14168;
  assign n14170 = ~n13889 & ~n14169;
  assign n14171 = ~n13893 & ~n13897;
  assign n14172 = ~n14170 & ~n14171;
  assign n14173 = ~n13870 & ~n13874;
  assign n14174 = ~n13873 & n14173;
  assign n14175 = ~n13869 & n14174;
  assign n14176 = ~n13867 & ~n14175;
  assign n14177 = ~n13871 & ~n13875;
  assign n14178 = ~n14176 & ~n14177;
  assign n14179 = ~n14172 & n14178;
  assign n14180 = n14172 & ~n14178;
  assign n14181 = ~n14179 & ~n14180;
  assign n14182 = ~n14166 & ~n14181;
  assign n14183 = ~n14165 & ~n14179;
  assign n14184 = ~n14180 & n14183;
  assign n14185 = ~n14162 & n14184;
  assign n14186 = ~n14182 & ~n14185;
  assign n14187 = ~n13829 & ~n13851;
  assign n14188 = ~n13807 & ~n14187;
  assign n14189 = ~n13828 & ~n13850;
  assign n14190 = ~n13847 & n14189;
  assign n14191 = ~n13825 & n14190;
  assign n14192 = ~n14188 & ~n14191;
  assign n14193 = ~n13838 & ~n13842;
  assign n14194 = ~n13841 & n14193;
  assign n14195 = ~n13837 & n14194;
  assign n14196 = ~n13835 & ~n14195;
  assign n14197 = ~n13839 & ~n13843;
  assign n14198 = ~n14196 & ~n14197;
  assign n14199 = ~n13816 & ~n13820;
  assign n14200 = ~n13819 & n14199;
  assign n14201 = ~n13815 & n14200;
  assign n14202 = ~n13813 & ~n14201;
  assign n14203 = ~n13817 & ~n13821;
  assign n14204 = ~n14202 & ~n14203;
  assign n14205 = ~n14198 & n14204;
  assign n14206 = n14198 & ~n14204;
  assign n14207 = ~n14205 & ~n14206;
  assign n14208 = ~n14192 & ~n14207;
  assign n14209 = ~n14191 & ~n14205;
  assign n14210 = ~n14206 & n14209;
  assign n14211 = ~n14188 & n14210;
  assign n14212 = ~n14208 & ~n14211;
  assign n14213 = ~n14186 & n14212;
  assign n14214 = n14186 & ~n14212;
  assign n14215 = ~n14213 & ~n14214;
  assign n14216 = ~n14160 & ~n14215;
  assign n14217 = n14160 & n14215;
  assign n14218 = ~n14216 & ~n14217;
  assign n14219 = ~n13739 & ~n13793;
  assign n14220 = ~n13685 & ~n14219;
  assign n14221 = n13739 & n13793;
  assign n14222 = ~n14220 & ~n14221;
  assign n14223 = ~n13765 & ~n13787;
  assign n14224 = ~n13743 & ~n14223;
  assign n14225 = ~n13764 & ~n13786;
  assign n14226 = ~n13783 & n14225;
  assign n14227 = ~n13761 & n14226;
  assign n14228 = ~n14224 & ~n14227;
  assign n14229 = ~n13774 & ~n13778;
  assign n14230 = ~n13777 & n14229;
  assign n14231 = ~n13773 & n14230;
  assign n14232 = ~n13771 & ~n14231;
  assign n14233 = ~n13775 & ~n13779;
  assign n14234 = ~n14232 & ~n14233;
  assign n14235 = ~n13752 & ~n13756;
  assign n14236 = ~n13755 & n14235;
  assign n14237 = ~n13751 & n14236;
  assign n14238 = ~n13749 & ~n14237;
  assign n14239 = ~n13753 & ~n13757;
  assign n14240 = ~n14238 & ~n14239;
  assign n14241 = ~n14234 & n14240;
  assign n14242 = n14234 & ~n14240;
  assign n14243 = ~n14241 & ~n14242;
  assign n14244 = ~n14228 & ~n14243;
  assign n14245 = ~n14227 & ~n14241;
  assign n14246 = ~n14242 & n14245;
  assign n14247 = ~n14224 & n14246;
  assign n14248 = ~n14244 & ~n14247;
  assign n14249 = ~n13711 & ~n13733;
  assign n14250 = ~n13689 & ~n14249;
  assign n14251 = ~n13710 & ~n13732;
  assign n14252 = ~n13729 & n14251;
  assign n14253 = ~n13707 & n14252;
  assign n14254 = ~n14250 & ~n14253;
  assign n14255 = ~n13720 & ~n13724;
  assign n14256 = ~n13723 & n14255;
  assign n14257 = ~n13719 & n14256;
  assign n14258 = ~n13717 & ~n14257;
  assign n14259 = ~n13721 & ~n13725;
  assign n14260 = ~n14258 & ~n14259;
  assign n14261 = ~n13698 & ~n13702;
  assign n14262 = ~n13701 & n14261;
  assign n14263 = ~n13697 & n14262;
  assign n14264 = ~n13695 & ~n14263;
  assign n14265 = ~n13699 & ~n13703;
  assign n14266 = ~n14264 & ~n14265;
  assign n14267 = ~n14260 & n14266;
  assign n14268 = n14260 & ~n14266;
  assign n14269 = ~n14267 & ~n14268;
  assign n14270 = ~n14254 & ~n14269;
  assign n14271 = ~n14253 & ~n14267;
  assign n14272 = ~n14268 & n14271;
  assign n14273 = ~n14250 & n14272;
  assign n14274 = ~n14270 & ~n14273;
  assign n14275 = ~n14248 & n14274;
  assign n14276 = n14248 & ~n14274;
  assign n14277 = ~n14275 & ~n14276;
  assign n14278 = ~n14222 & ~n14277;
  assign n14279 = n14222 & n14277;
  assign n14280 = ~n14278 & ~n14279;
  assign n14281 = ~n14218 & n14280;
  assign n14282 = n14218 & ~n14280;
  assign n14283 = ~n14281 & ~n14282;
  assign n14284 = ~n14156 & ~n14283;
  assign n14285 = n14156 & n14283;
  assign n14286 = ~n14284 & ~n14285;
  assign n14287 = ~n14152 & ~n14286;
  assign n14288 = ~n13928 & ~n14287;
  assign n14289 = ~n14150 & n14286;
  assign n14290 = ~n14151 & n14289;
  assign n14291 = ~n14288 & ~n14290;
  assign n14292 = ~n14066 & ~n14146;
  assign n14293 = ~n13932 & ~n14292;
  assign n14294 = n14066 & n14146;
  assign n14295 = ~n14293 & ~n14294;
  assign n14296 = ~n14113 & ~n14139;
  assign n14297 = ~n14071 & ~n14296;
  assign n14298 = ~n14109 & n14139;
  assign n14299 = ~n14112 & n14298;
  assign n14300 = ~n14297 & ~n14299;
  assign n14301 = ~n14124 & ~n14130;
  assign n14302 = ~n14129 & n14301;
  assign n14303 = ~n14123 & n14302;
  assign n14304 = ~n14119 & ~n14303;
  assign n14305 = ~n14125 & ~n14131;
  assign n14306 = ~n14304 & ~n14305;
  assign n14307 = n14103 & ~n14106;
  assign n14308 = ~n14076 & ~n14307;
  assign n14309 = ~n14097 & ~n14103;
  assign n14310 = ~n14094 & n14309;
  assign n14311 = ~n14308 & ~n14310;
  assign n14312 = ~n13302 & ~n14087;
  assign n14313 = ~n14089 & n14312;
  assign n14314 = ~n14086 & n14313;
  assign n14315 = ~n14082 & ~n14314;
  assign n14316 = ~n14088 & ~n14090;
  assign n14317 = ~n14315 & ~n14316;
  assign n14318 = ~n14311 & n14317;
  assign n14319 = ~n14310 & ~n14317;
  assign n14320 = ~n14308 & n14319;
  assign n14321 = ~n14318 & ~n14320;
  assign n14322 = ~n14306 & ~n14321;
  assign n14323 = n14306 & ~n14320;
  assign n14324 = ~n14318 & n14323;
  assign n14325 = ~n14322 & ~n14324;
  assign n14326 = ~n14300 & n14325;
  assign n14327 = n14300 & ~n14325;
  assign n14328 = ~n14326 & ~n14327;
  assign n14329 = ~n13998 & ~n14060;
  assign n14330 = ~n13936 & ~n14329;
  assign n14331 = n13998 & n14060;
  assign n14332 = ~n14330 & ~n14331;
  assign n14333 = ~n14028 & ~n14054;
  assign n14334 = ~n14002 & ~n14333;
  assign n14335 = ~n14027 & ~n14053;
  assign n14336 = ~n14050 & n14335;
  assign n14337 = ~n14024 & n14336;
  assign n14338 = ~n14334 & ~n14337;
  assign n14339 = ~n14013 & ~n14019;
  assign n14340 = ~n14018 & n14339;
  assign n14341 = ~n14012 & n14340;
  assign n14342 = ~n14008 & ~n14341;
  assign n14343 = ~n14014 & ~n14020;
  assign n14344 = ~n14342 & ~n14343;
  assign n14345 = ~n14039 & ~n14045;
  assign n14346 = ~n14044 & n14345;
  assign n14347 = ~n14038 & n14346;
  assign n14348 = ~n14034 & ~n14347;
  assign n14349 = ~n14040 & ~n14046;
  assign n14350 = ~n14348 & ~n14349;
  assign n14351 = ~n14344 & n14350;
  assign n14352 = n14344 & ~n14350;
  assign n14353 = ~n14351 & ~n14352;
  assign n14354 = ~n14338 & ~n14353;
  assign n14355 = ~n14337 & ~n14351;
  assign n14356 = ~n14352 & n14355;
  assign n14357 = ~n14334 & n14356;
  assign n14358 = ~n14354 & ~n14357;
  assign n14359 = ~n13966 & ~n13992;
  assign n14360 = ~n13940 & ~n14359;
  assign n14361 = ~n13965 & ~n13991;
  assign n14362 = ~n13988 & n14361;
  assign n14363 = ~n13962 & n14362;
  assign n14364 = ~n14360 & ~n14363;
  assign n14365 = ~n13951 & ~n13957;
  assign n14366 = ~n13956 & n14365;
  assign n14367 = ~n13950 & n14366;
  assign n14368 = ~n13946 & ~n14367;
  assign n14369 = ~n13952 & ~n13958;
  assign n14370 = ~n14368 & ~n14369;
  assign n14371 = ~n13977 & ~n13983;
  assign n14372 = ~n13982 & n14371;
  assign n14373 = ~n13976 & n14372;
  assign n14374 = ~n13972 & ~n14373;
  assign n14375 = ~n13978 & ~n13984;
  assign n14376 = ~n14374 & ~n14375;
  assign n14377 = ~n14370 & n14376;
  assign n14378 = n14370 & ~n14376;
  assign n14379 = ~n14377 & ~n14378;
  assign n14380 = ~n14364 & ~n14379;
  assign n14381 = ~n14363 & ~n14377;
  assign n14382 = ~n14378 & n14381;
  assign n14383 = ~n14360 & n14382;
  assign n14384 = ~n14380 & ~n14383;
  assign n14385 = ~n14358 & n14384;
  assign n14386 = n14358 & ~n14384;
  assign n14387 = ~n14385 & ~n14386;
  assign n14388 = ~n14332 & ~n14387;
  assign n14389 = n14332 & n14387;
  assign n14390 = ~n14388 & ~n14389;
  assign n14391 = ~n14328 & n14390;
  assign n14392 = n14328 & ~n14390;
  assign n14393 = ~n14391 & ~n14392;
  assign n14394 = ~n14295 & ~n14393;
  assign n14395 = n14295 & n14393;
  assign n14396 = ~n14394 & ~n14395;
  assign n14397 = ~n14218 & ~n14280;
  assign n14398 = ~n14156 & ~n14397;
  assign n14399 = n14218 & n14280;
  assign n14400 = ~n14398 & ~n14399;
  assign n14401 = ~n14248 & ~n14274;
  assign n14402 = ~n14222 & ~n14401;
  assign n14403 = ~n14247 & ~n14273;
  assign n14404 = ~n14270 & n14403;
  assign n14405 = ~n14244 & n14404;
  assign n14406 = ~n14402 & ~n14405;
  assign n14407 = ~n14233 & ~n14239;
  assign n14408 = ~n14238 & n14407;
  assign n14409 = ~n14232 & n14408;
  assign n14410 = ~n14228 & ~n14409;
  assign n14411 = ~n14234 & ~n14240;
  assign n14412 = ~n14410 & ~n14411;
  assign n14413 = ~n14259 & ~n14265;
  assign n14414 = ~n14264 & n14413;
  assign n14415 = ~n14258 & n14414;
  assign n14416 = ~n14254 & ~n14415;
  assign n14417 = ~n14260 & ~n14266;
  assign n14418 = ~n14416 & ~n14417;
  assign n14419 = ~n14412 & n14418;
  assign n14420 = n14412 & ~n14418;
  assign n14421 = ~n14419 & ~n14420;
  assign n14422 = ~n14406 & ~n14421;
  assign n14423 = ~n14405 & ~n14419;
  assign n14424 = ~n14420 & n14423;
  assign n14425 = ~n14402 & n14424;
  assign n14426 = ~n14422 & ~n14425;
  assign n14427 = ~n14186 & ~n14212;
  assign n14428 = ~n14160 & ~n14427;
  assign n14429 = ~n14185 & ~n14211;
  assign n14430 = ~n14208 & n14429;
  assign n14431 = ~n14182 & n14430;
  assign n14432 = ~n14428 & ~n14431;
  assign n14433 = ~n14171 & ~n14177;
  assign n14434 = ~n14176 & n14433;
  assign n14435 = ~n14170 & n14434;
  assign n14436 = ~n14166 & ~n14435;
  assign n14437 = ~n14172 & ~n14178;
  assign n14438 = ~n14436 & ~n14437;
  assign n14439 = ~n14197 & ~n14203;
  assign n14440 = ~n14202 & n14439;
  assign n14441 = ~n14196 & n14440;
  assign n14442 = ~n14192 & ~n14441;
  assign n14443 = ~n14198 & ~n14204;
  assign n14444 = ~n14442 & ~n14443;
  assign n14445 = ~n14438 & n14444;
  assign n14446 = n14438 & ~n14444;
  assign n14447 = ~n14445 & ~n14446;
  assign n14448 = ~n14432 & ~n14447;
  assign n14449 = ~n14431 & ~n14445;
  assign n14450 = ~n14446 & n14449;
  assign n14451 = ~n14428 & n14450;
  assign n14452 = ~n14448 & ~n14451;
  assign n14453 = ~n14426 & n14452;
  assign n14454 = n14426 & ~n14452;
  assign n14455 = ~n14453 & ~n14454;
  assign n14456 = ~n14400 & ~n14455;
  assign n14457 = n14400 & n14455;
  assign n14458 = ~n14456 & ~n14457;
  assign n14459 = ~n14396 & ~n14458;
  assign n14460 = ~n14291 & ~n14459;
  assign n14461 = ~n14394 & n14458;
  assign n14462 = ~n14395 & n14461;
  assign n14463 = ~n14460 & ~n14462;
  assign n14464 = ~n14328 & ~n14390;
  assign n14465 = ~n14295 & ~n14464;
  assign n14466 = n14328 & n14390;
  assign n14467 = ~n14465 & ~n14466;
  assign n14468 = ~n14300 & ~n14324;
  assign n14469 = ~n14322 & ~n14468;
  assign n14470 = ~n14311 & ~n14317;
  assign n14471 = ~n14469 & n14470;
  assign n14472 = ~n14322 & ~n14470;
  assign n14473 = ~n14468 & n14472;
  assign n14474 = ~n14471 & ~n14473;
  assign n14475 = ~n14358 & ~n14384;
  assign n14476 = ~n14332 & ~n14475;
  assign n14477 = ~n14357 & ~n14383;
  assign n14478 = ~n14380 & n14477;
  assign n14479 = ~n14354 & n14478;
  assign n14480 = ~n14476 & ~n14479;
  assign n14481 = ~n14369 & ~n14375;
  assign n14482 = ~n14374 & n14481;
  assign n14483 = ~n14368 & n14482;
  assign n14484 = ~n14364 & ~n14483;
  assign n14485 = ~n14370 & ~n14376;
  assign n14486 = ~n14484 & ~n14485;
  assign n14487 = ~n14343 & ~n14349;
  assign n14488 = ~n14348 & n14487;
  assign n14489 = ~n14342 & n14488;
  assign n14490 = ~n14338 & ~n14489;
  assign n14491 = ~n14344 & ~n14350;
  assign n14492 = ~n14490 & ~n14491;
  assign n14493 = ~n14486 & n14492;
  assign n14494 = n14486 & ~n14492;
  assign n14495 = ~n14493 & ~n14494;
  assign n14496 = ~n14480 & ~n14495;
  assign n14497 = ~n14479 & ~n14493;
  assign n14498 = ~n14494 & n14497;
  assign n14499 = ~n14476 & n14498;
  assign n14500 = ~n14496 & ~n14499;
  assign n14501 = ~n14474 & ~n14500;
  assign n14502 = ~n14473 & ~n14499;
  assign n14503 = ~n14471 & n14502;
  assign n14504 = ~n14496 & n14503;
  assign n14505 = ~n14501 & ~n14504;
  assign n14506 = ~n14467 & n14505;
  assign n14507 = n14467 & ~n14505;
  assign n14508 = ~n14506 & ~n14507;
  assign n14509 = ~n14426 & ~n14452;
  assign n14510 = ~n14400 & ~n14509;
  assign n14511 = ~n14425 & ~n14451;
  assign n14512 = ~n14448 & n14511;
  assign n14513 = ~n14422 & n14512;
  assign n14514 = ~n14510 & ~n14513;
  assign n14515 = ~n14437 & ~n14443;
  assign n14516 = ~n14442 & n14515;
  assign n14517 = ~n14436 & n14516;
  assign n14518 = ~n14432 & ~n14517;
  assign n14519 = ~n14438 & ~n14444;
  assign n14520 = ~n14518 & ~n14519;
  assign n14521 = ~n14411 & ~n14417;
  assign n14522 = ~n14416 & n14521;
  assign n14523 = ~n14410 & n14522;
  assign n14524 = ~n14406 & ~n14523;
  assign n14525 = ~n14412 & ~n14418;
  assign n14526 = ~n14524 & ~n14525;
  assign n14527 = ~n14520 & n14526;
  assign n14528 = n14520 & ~n14526;
  assign n14529 = ~n14527 & ~n14528;
  assign n14530 = ~n14514 & ~n14529;
  assign n14531 = ~n14513 & ~n14527;
  assign n14532 = ~n14528 & n14531;
  assign n14533 = ~n14510 & n14532;
  assign n14534 = ~n14530 & ~n14533;
  assign n14535 = ~n14508 & ~n14534;
  assign n14536 = ~n14463 & ~n14535;
  assign n14537 = ~n14506 & n14534;
  assign n14538 = ~n14507 & n14537;
  assign n14539 = ~n14536 & ~n14538;
  assign n14540 = ~n14467 & ~n14501;
  assign n14541 = ~n14504 & ~n14540;
  assign n14542 = ~n14485 & ~n14491;
  assign n14543 = ~n14490 & n14542;
  assign n14544 = ~n14484 & n14543;
  assign n14545 = ~n14480 & ~n14544;
  assign n14546 = ~n14486 & ~n14492;
  assign n14547 = ~n14471 & ~n14546;
  assign n14548 = ~n14545 & n14547;
  assign n14549 = ~n14545 & ~n14546;
  assign n14550 = n14471 & ~n14549;
  assign n14551 = ~n14548 & ~n14550;
  assign n14552 = ~n14541 & n14551;
  assign n14553 = ~n14504 & ~n14551;
  assign n14554 = ~n14540 & n14553;
  assign n14555 = ~n14552 & ~n14554;
  assign n14556 = ~n14519 & ~n14525;
  assign n14557 = ~n14524 & n14556;
  assign n14558 = ~n14518 & n14557;
  assign n14559 = ~n14514 & ~n14558;
  assign n14560 = ~n14520 & ~n14526;
  assign n14561 = ~n14559 & ~n14560;
  assign n14562 = ~n14555 & n14561;
  assign n14563 = ~n14539 & ~n14562;
  assign n14564 = ~n14554 & ~n14561;
  assign n14565 = ~n14552 & n14564;
  assign n14566 = ~n14563 & ~n14565;
  assign n14567 = ~n14541 & ~n14548;
  assign n14568 = ~n14550 & ~n14567;
  assign n14569 = ~n14566 & n14568;
  assign n14570 = ~n14565 & ~n14568;
  assign n14571 = ~n14563 & n14570;
  assign n14572 = ~n14569 & ~n14571;
  assign n14573 = ~n14555 & ~n14561;
  assign n14574 = ~n14554 & n14561;
  assign n14575 = ~n14552 & n14574;
  assign n14576 = ~n14538 & ~n14575;
  assign n14577 = ~n14536 & n14576;
  assign n14578 = ~n14573 & n14577;
  assign n14579 = ~n14573 & ~n14575;
  assign n14580 = ~n14539 & ~n14579;
  assign n14581 = ~n14508 & n14534;
  assign n14582 = ~n14506 & ~n14534;
  assign n14583 = ~n14507 & n14582;
  assign n14584 = ~n14581 & ~n14583;
  assign n14585 = n14463 & n14584;
  assign n14586 = ~n14463 & ~n14584;
  assign n14587 = ~n14394 & ~n14458;
  assign n14588 = ~n14395 & n14587;
  assign n14589 = ~n14396 & n14458;
  assign n14590 = ~n14588 & ~n14589;
  assign n14591 = n14291 & n14590;
  assign n14592 = ~n14291 & ~n14590;
  assign n14593 = ~n14152 & n14286;
  assign n14594 = ~n14150 & ~n14286;
  assign n14595 = ~n14151 & n14594;
  assign n14596 = ~n14593 & ~n14595;
  assign n14597 = n13928 & n14596;
  assign n14598 = ~n13928 & ~n14596;
  assign n14599 = ~n13675 & ~n13923;
  assign n14600 = ~n13676 & n14599;
  assign n14601 = ~n13677 & n13923;
  assign n14602 = ~n14600 & ~n14601;
  assign n14603 = n13275 & n14602;
  assign n14604 = ~n13275 & ~n14602;
  assign n14605 = ~n12736 & n13270;
  assign n14606 = ~n12734 & ~n13270;
  assign n14607 = ~n12735 & n14606;
  assign n14608 = ~n14605 & ~n14607;
  assign n14609 = n11871 & n14608;
  assign n14610 = ~n11871 & ~n14608;
  assign n14611 = ~n11168 & ~n11866;
  assign n14612 = ~n11169 & n14611;
  assign n14613 = ~n11170 & n11866;
  assign n14614 = ~n14612 & ~n14613;
  assign n14615 = ~n10047 & ~n14614;
  assign n14616 = ~n10032 & ~n10033;
  assign n14617 = ~n10034 & n14616;
  assign n14618 = n10032 & ~n10035;
  assign n14619 = ~n14617 & ~n14618;
  assign n14620 = A1000  & ~n14619;
  assign n14621 = ~n14615 & n14620;
  assign n14622 = n10047 & n14614;
  assign n14623 = n10036 & ~n10041;
  assign n14624 = ~n10029 & n14623;
  assign n14625 = ~n10036 & ~n10045;
  assign n14626 = ~n14624 & ~n14625;
  assign n14627 = n4472 & ~n14626;
  assign n14628 = ~n10043 & ~n10046;
  assign n14629 = ~n4472 & ~n14628;
  assign n14630 = ~n14627 & ~n14629;
  assign n14631 = ~n14622 & ~n14630;
  assign n14632 = n14621 & n14631;
  assign n14633 = ~n14610 & n14632;
  assign n14634 = ~n14609 & n14633;
  assign n14635 = ~n14604 & n14634;
  assign n14636 = ~n14603 & n14635;
  assign n14637 = ~n14598 & n14636;
  assign n14638 = ~n14597 & n14637;
  assign n14639 = ~n14592 & n14638;
  assign n14640 = ~n14591 & n14639;
  assign n14641 = ~n14586 & n14640;
  assign n14642 = ~n14585 & n14641;
  assign n14643 = ~n14580 & n14642;
  assign n14644 = ~n14578 & n14643;
  assign n14645 = n14572 & n14644;
  assign n14646 = ~n14572 & ~n14644;
  assign n14647 = ~n14645 & ~n14646;
  assign n14648 = ~n14578 & ~n14580;
  assign n14649 = ~n14642 & ~n14648;
  assign n14650 = ~n14585 & ~n14586;
  assign n14651 = ~n14640 & ~n14650;
  assign n14652 = ~n14591 & ~n14592;
  assign n14653 = ~n14638 & ~n14652;
  assign n14654 = ~n14609 & ~n14610;
  assign n14655 = ~n14632 & ~n14654;
  assign n14656 = ~n14615 & ~n14622;
  assign n14657 = n14620 & ~n14630;
  assign n14658 = ~n14656 & ~n14657;
  assign n14659 = ~n14632 & ~n14658;
  assign n14660 = n14620 & ~n14627;
  assign n14661 = ~n14629 & n14660;
  assign n14662 = ~n14620 & ~n14630;
  assign n14663 = ~n14661 & ~n14662;
  assign n14664 = ~n14659 & n14663;
  assign n14665 = ~n14634 & ~n14664;
  assign n14666 = ~n14655 & n14665;
  assign n14667 = ~n14603 & ~n14604;
  assign n14668 = ~n14634 & ~n14667;
  assign n14669 = ~n14636 & ~n14668;
  assign n14670 = ~n14666 & ~n14669;
  assign n14671 = ~n14597 & ~n14598;
  assign n14672 = ~n14636 & ~n14671;
  assign n14673 = ~n14638 & ~n14672;
  assign n14674 = ~n14670 & n14673;
  assign n14675 = ~n14640 & n14674;
  assign n14676 = ~n14653 & n14675;
  assign n14677 = ~n14642 & n14676;
  assign n14678 = ~n14651 & n14677;
  assign n14679 = ~n14644 & n14678;
  assign n14680 = ~n14649 & n14679;
  assign n14681 = ~n14647 & n14680;
  assign n14682 = ~n14572 & n14644;
  assign n14683 = ~n14566 & ~n14568;
  assign n14684 = ~n14682 & n14683;
  assign n14685 = n14644 & ~n14683;
  assign n14686 = ~n14572 & n14685;
  assign n14687 = ~n14568 & n14640;
  assign n14688 = n14650 & n14687;
  assign n14689 = ~n14580 & n14688;
  assign n14690 = ~n14578 & n14689;
  assign n14691 = ~n14566 & n14690;
  assign n14692 = ~n14572 & n14691;
  assign n14693 = ~n14686 & ~n14692;
  assign n14694 = ~n14684 & n14693;
  assign n14695 = ~n14681 & n14694;
  assign n14696 = ~n14642 & ~n14651;
  assign n14697 = ~n14634 & ~n14655;
  assign n14698 = n14664 & ~n14697;
  assign n14699 = ~n14666 & ~n14698;
  assign n14700 = n14659 & ~n14663;
  assign n14701 = A1000  & ~n14617;
  assign n14702 = ~n14618 & n14701;
  assign n14703 = ~A1000  & ~n14619;
  assign n14704 = ~n14702 & ~n14703;
  assign n14705 = ~n14664 & n14704;
  assign n14706 = ~n14700 & n14705;
  assign n14707 = n14659 & ~n14706;
  assign n14708 = ~n14664 & ~n14700;
  assign n14709 = ~n14704 & ~n14708;
  assign n14710 = ~n14707 & ~n14709;
  assign n14711 = ~n14699 & n14710;
  assign n14712 = n14697 & ~n14711;
  assign n14713 = n14699 & ~n14710;
  assign n14714 = ~n14712 & ~n14713;
  assign n14715 = ~n14666 & ~n14714;
  assign n14716 = ~n14636 & n14666;
  assign n14717 = ~n14668 & n14716;
  assign n14718 = n14670 & ~n14673;
  assign n14719 = ~n14674 & ~n14718;
  assign n14720 = ~n14717 & ~n14719;
  assign n14721 = ~n14715 & n14720;
  assign n14722 = n14673 & ~n14721;
  assign n14723 = ~n14715 & ~n14717;
  assign n14724 = n14719 & ~n14723;
  assign n14725 = ~n14722 & ~n14724;
  assign n14726 = n14674 & ~n14725;
  assign n14727 = ~n14640 & ~n14653;
  assign n14728 = ~n14674 & n14727;
  assign n14729 = ~n14676 & ~n14696;
  assign n14730 = ~n14678 & ~n14729;
  assign n14731 = ~n14728 & ~n14730;
  assign n14732 = ~n14726 & n14731;
  assign n14733 = n14696 & ~n14732;
  assign n14734 = ~n14726 & ~n14728;
  assign n14735 = n14730 & ~n14734;
  assign n14736 = ~n14733 & ~n14735;
  assign n14737 = n14678 & ~n14680;
  assign n14738 = ~n14736 & n14737;
  assign n14739 = n14680 & ~n14733;
  assign n14740 = ~n14735 & n14739;
  assign n14741 = ~n14644 & ~n14649;
  assign n14742 = ~n14740 & n14741;
  assign n14743 = ~n14738 & ~n14742;
  assign n14744 = n14680 & ~n14681;
  assign n14745 = ~n14743 & n14744;
  assign n14746 = n14681 & ~n14738;
  assign n14747 = ~n14742 & n14746;
  assign n14748 = ~n14647 & ~n14747;
  assign n14749 = ~n14681 & ~n14748;
  assign n14750 = ~n14745 & n14749;
  assign n14751 = n14680 & ~n14686;
  assign n14752 = ~n14684 & n14751;
  assign n14753 = ~n14647 & n14752;
  assign n14754 = ~n14684 & ~n14686;
  assign n14755 = ~n14681 & n14754;
  assign n14756 = n14692 & ~n14755;
  assign n14757 = ~n14695 & ~n14756;
  assign n14758 = ~n14753 & ~n14757;
  assign n14759 = ~n14750 & n14758;
  assign maj = ~n14695 | n14759;
endmodule


